VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO alu_32_bit
  CLASS BLOCK ;
  FOREIGN alu_32_bit ;
  ORIGIN 0.000 0.000 ;
  SIZE 434.090 BY 444.810 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 430.090 435.240 434.090 435.840 ;
    END
  END A[0]
  PIN A[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 430.090 418.240 434.090 418.840 ;
    END
  END A[10]
  PIN A[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END A[11]
  PIN A[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END A[12]
  PIN A[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END A[13]
  PIN A[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 430.090 292.440 434.090 293.040 ;
    END
  END A[14]
  PIN A[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 430.090 149.640 434.090 150.240 ;
    END
  END A[15]
  PIN A[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END A[16]
  PIN A[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 430.090 57.840 434.090 58.440 ;
    END
  END A[17]
  PIN A[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END A[18]
  PIN A[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END A[19]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END A[1]
  PIN A[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END A[20]
  PIN A[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 289.890 440.810 290.170 444.810 ;
    END
  END A[21]
  PIN A[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 103.130 440.810 103.410 444.810 ;
    END
  END A[22]
  PIN A[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 119.230 440.810 119.510 444.810 ;
    END
  END A[23]
  PIN A[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 430.090 238.040 434.090 238.640 ;
    END
  END A[24]
  PIN A[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END A[25]
  PIN A[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 430.090 397.840 434.090 398.440 ;
    END
  END A[26]
  PIN A[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END A[27]
  PIN A[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 430.090 326.440 434.090 327.040 ;
    END
  END A[28]
  PIN A[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END A[29]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END A[2]
  PIN A[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END A[30]
  PIN A[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 270.570 440.810 270.850 444.810 ;
    END
  END A[31]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 430.090 221.040 434.090 221.640 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 154.650 440.810 154.930 444.810 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 170.750 440.810 171.030 444.810 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 430.090 380.840 434.090 381.440 ;
    END
  END A[9]
  PIN B[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 430.090 95.240 434.090 95.840 ;
    END
  END B[0]
  PIN B[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 254.470 440.810 254.750 444.810 ;
    END
  END B[10]
  PIN B[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 430.090 129.240 434.090 129.840 ;
    END
  END B[11]
  PIN B[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 186.850 440.810 187.130 444.810 ;
    END
  END B[12]
  PIN B[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 322.090 440.810 322.370 444.810 ;
    END
  END B[13]
  PIN B[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END B[14]
  PIN B[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END B[15]
  PIN B[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 430.090 23.840 434.090 24.440 ;
    END
  END B[16]
  PIN B[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 430.090 363.840 434.090 364.440 ;
    END
  END B[17]
  PIN B[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 430.090 183.640 434.090 184.240 ;
    END
  END B[18]
  PIN B[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 222.270 440.810 222.550 444.810 ;
    END
  END B[19]
  PIN B[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 357.510 440.810 357.790 444.810 ;
    END
  END B[1]
  PIN B[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 430.090 3.440 434.090 4.040 ;
    END
  END B[20]
  PIN B[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 430.090 346.840 434.090 347.440 ;
    END
  END B[21]
  PIN B[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 409.030 440.810 409.310 444.810 ;
    END
  END B[22]
  PIN B[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 238.370 440.810 238.650 444.810 ;
    END
  END B[23]
  PIN B[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END B[24]
  PIN B[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 430.090 78.240 434.090 78.840 ;
    END
  END B[25]
  PIN B[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END B[26]
  PIN B[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END B[27]
  PIN B[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END B[28]
  PIN B[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END B[29]
  PIN B[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 135.330 440.810 135.610 444.810 ;
    END
  END B[2]
  PIN B[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 373.610 440.810 373.890 444.810 ;
    END
  END B[30]
  PIN B[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END B[31]
  PIN B[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END B[3]
  PIN B[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END B[4]
  PIN B[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END B[5]
  PIN B[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END B[6]
  PIN B[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 430.090 112.240 434.090 112.840 ;
    END
  END B[7]
  PIN B[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END B[8]
  PIN B[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END B[9]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 432.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 428.500 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 428.500 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 428.500 337.990 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 432.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 432.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 428.500 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 428.500 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 428.500 334.690 ;
    END
  END VPWR
  PIN control[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END control[0]
  PIN control[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 51.610 440.810 51.890 444.810 ;
    END
  END control[1]
  PIN control[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 430.090 166.640 434.090 167.240 ;
    END
  END control[2]
  PIN control[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END control[3]
  PIN result[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END result[0]
  PIN result[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 430.090 309.440 434.090 310.040 ;
    END
  END result[10]
  PIN result[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 67.710 440.810 67.990 444.810 ;
    END
  END result[11]
  PIN result[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END result[12]
  PIN result[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END result[13]
  PIN result[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END result[14]
  PIN result[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END result[15]
  PIN result[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END result[16]
  PIN result[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 202.950 440.810 203.230 444.810 ;
    END
  END result[17]
  PIN result[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END result[18]
  PIN result[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 440.810 0.370 444.810 ;
    END
  END result[19]
  PIN result[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END result[1]
  PIN result[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END result[20]
  PIN result[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 389.710 440.810 389.990 444.810 ;
    END
  END result[21]
  PIN result[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 305.990 440.810 306.270 444.810 ;
    END
  END result[22]
  PIN result[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END result[23]
  PIN result[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 425.130 440.810 425.410 444.810 ;
    END
  END result[24]
  PIN result[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 430.090 40.840 434.090 41.440 ;
    END
  END result[25]
  PIN result[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 16.190 440.810 16.470 444.810 ;
    END
  END result[26]
  PIN result[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 430.090 255.040 434.090 255.640 ;
    END
  END result[27]
  PIN result[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END result[28]
  PIN result[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END result[29]
  PIN result[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END result[2]
  PIN result[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 430.090 272.040 434.090 272.640 ;
    END
  END result[30]
  PIN result[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END result[31]
  PIN result[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END result[3]
  PIN result[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 341.410 440.810 341.690 444.810 ;
    END
  END result[4]
  PIN result[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 35.510 440.810 35.790 444.810 ;
    END
  END result[5]
  PIN result[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 87.030 440.810 87.310 444.810 ;
    END
  END result[6]
  PIN result[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END result[7]
  PIN result[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END result[8]
  PIN result[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END result[9]
  PIN zero_flag
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 430.090 200.640 434.090 201.240 ;
    END
  END zero_flag
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 428.260 432.565 ;
      LAYER met1 ;
        RECT 0.070 10.640 428.650 432.720 ;
      LAYER met2 ;
        RECT 0.650 440.530 15.910 440.810 ;
        RECT 16.750 440.530 35.230 440.810 ;
        RECT 36.070 440.530 51.330 440.810 ;
        RECT 52.170 440.530 67.430 440.810 ;
        RECT 68.270 440.530 86.750 440.810 ;
        RECT 87.590 440.530 102.850 440.810 ;
        RECT 103.690 440.530 118.950 440.810 ;
        RECT 119.790 440.530 135.050 440.810 ;
        RECT 135.890 440.530 154.370 440.810 ;
        RECT 155.210 440.530 170.470 440.810 ;
        RECT 171.310 440.530 186.570 440.810 ;
        RECT 187.410 440.530 202.670 440.810 ;
        RECT 203.510 440.530 221.990 440.810 ;
        RECT 222.830 440.530 238.090 440.810 ;
        RECT 238.930 440.530 254.190 440.810 ;
        RECT 255.030 440.530 270.290 440.810 ;
        RECT 271.130 440.530 289.610 440.810 ;
        RECT 290.450 440.530 305.710 440.810 ;
        RECT 306.550 440.530 321.810 440.810 ;
        RECT 322.650 440.530 341.130 440.810 ;
        RECT 341.970 440.530 357.230 440.810 ;
        RECT 358.070 440.530 373.330 440.810 ;
        RECT 374.170 440.530 389.430 440.810 ;
        RECT 390.270 440.530 408.750 440.810 ;
        RECT 409.590 440.530 424.850 440.810 ;
        RECT 425.690 440.530 428.630 440.810 ;
        RECT 0.100 4.280 428.630 440.530 ;
        RECT 0.650 3.555 15.910 4.280 ;
        RECT 16.750 3.555 32.010 4.280 ;
        RECT 32.850 3.555 48.110 4.280 ;
        RECT 48.950 3.555 67.430 4.280 ;
        RECT 68.270 3.555 83.530 4.280 ;
        RECT 84.370 3.555 99.630 4.280 ;
        RECT 100.470 3.555 115.730 4.280 ;
        RECT 116.570 3.555 135.050 4.280 ;
        RECT 135.890 3.555 151.150 4.280 ;
        RECT 151.990 3.555 167.250 4.280 ;
        RECT 168.090 3.555 183.350 4.280 ;
        RECT 184.190 3.555 202.670 4.280 ;
        RECT 203.510 3.555 218.770 4.280 ;
        RECT 219.610 3.555 234.870 4.280 ;
        RECT 235.710 3.555 254.190 4.280 ;
        RECT 255.030 3.555 270.290 4.280 ;
        RECT 271.130 3.555 286.390 4.280 ;
        RECT 287.230 3.555 302.490 4.280 ;
        RECT 303.330 3.555 321.810 4.280 ;
        RECT 322.650 3.555 337.910 4.280 ;
        RECT 338.750 3.555 354.010 4.280 ;
        RECT 354.850 3.555 370.110 4.280 ;
        RECT 370.950 3.555 389.430 4.280 ;
        RECT 390.270 3.555 405.530 4.280 ;
        RECT 406.370 3.555 421.630 4.280 ;
        RECT 422.470 3.555 428.630 4.280 ;
      LAYER met3 ;
        RECT 3.990 434.840 429.690 435.705 ;
        RECT 3.990 429.440 430.090 434.840 ;
        RECT 4.400 428.040 430.090 429.440 ;
        RECT 3.990 419.240 430.090 428.040 ;
        RECT 3.990 417.840 429.690 419.240 ;
        RECT 3.990 412.440 430.090 417.840 ;
        RECT 4.400 411.040 430.090 412.440 ;
        RECT 3.990 398.840 430.090 411.040 ;
        RECT 3.990 397.440 429.690 398.840 ;
        RECT 3.990 392.040 430.090 397.440 ;
        RECT 4.400 390.640 430.090 392.040 ;
        RECT 3.990 381.840 430.090 390.640 ;
        RECT 3.990 380.440 429.690 381.840 ;
        RECT 3.990 375.040 430.090 380.440 ;
        RECT 4.400 373.640 430.090 375.040 ;
        RECT 3.990 364.840 430.090 373.640 ;
        RECT 3.990 363.440 429.690 364.840 ;
        RECT 3.990 358.040 430.090 363.440 ;
        RECT 4.400 356.640 430.090 358.040 ;
        RECT 3.990 347.840 430.090 356.640 ;
        RECT 3.990 346.440 429.690 347.840 ;
        RECT 3.990 341.040 430.090 346.440 ;
        RECT 4.400 339.640 430.090 341.040 ;
        RECT 3.990 327.440 430.090 339.640 ;
        RECT 3.990 326.040 429.690 327.440 ;
        RECT 3.990 320.640 430.090 326.040 ;
        RECT 4.400 319.240 430.090 320.640 ;
        RECT 3.990 310.440 430.090 319.240 ;
        RECT 3.990 309.040 429.690 310.440 ;
        RECT 3.990 303.640 430.090 309.040 ;
        RECT 4.400 302.240 430.090 303.640 ;
        RECT 3.990 293.440 430.090 302.240 ;
        RECT 3.990 292.040 429.690 293.440 ;
        RECT 3.990 286.640 430.090 292.040 ;
        RECT 4.400 285.240 430.090 286.640 ;
        RECT 3.990 273.040 430.090 285.240 ;
        RECT 3.990 271.640 429.690 273.040 ;
        RECT 3.990 269.640 430.090 271.640 ;
        RECT 4.400 268.240 430.090 269.640 ;
        RECT 3.990 256.040 430.090 268.240 ;
        RECT 3.990 254.640 429.690 256.040 ;
        RECT 3.990 249.240 430.090 254.640 ;
        RECT 4.400 247.840 430.090 249.240 ;
        RECT 3.990 239.040 430.090 247.840 ;
        RECT 3.990 237.640 429.690 239.040 ;
        RECT 3.990 232.240 430.090 237.640 ;
        RECT 4.400 230.840 430.090 232.240 ;
        RECT 3.990 222.040 430.090 230.840 ;
        RECT 3.990 220.640 429.690 222.040 ;
        RECT 3.990 215.240 430.090 220.640 ;
        RECT 4.400 213.840 430.090 215.240 ;
        RECT 3.990 201.640 430.090 213.840 ;
        RECT 3.990 200.240 429.690 201.640 ;
        RECT 3.990 194.840 430.090 200.240 ;
        RECT 4.400 193.440 430.090 194.840 ;
        RECT 3.990 184.640 430.090 193.440 ;
        RECT 3.990 183.240 429.690 184.640 ;
        RECT 3.990 177.840 430.090 183.240 ;
        RECT 4.400 176.440 430.090 177.840 ;
        RECT 3.990 167.640 430.090 176.440 ;
        RECT 3.990 166.240 429.690 167.640 ;
        RECT 3.990 160.840 430.090 166.240 ;
        RECT 4.400 159.440 430.090 160.840 ;
        RECT 3.990 150.640 430.090 159.440 ;
        RECT 3.990 149.240 429.690 150.640 ;
        RECT 3.990 143.840 430.090 149.240 ;
        RECT 4.400 142.440 430.090 143.840 ;
        RECT 3.990 130.240 430.090 142.440 ;
        RECT 3.990 128.840 429.690 130.240 ;
        RECT 3.990 123.440 430.090 128.840 ;
        RECT 4.400 122.040 430.090 123.440 ;
        RECT 3.990 113.240 430.090 122.040 ;
        RECT 3.990 111.840 429.690 113.240 ;
        RECT 3.990 106.440 430.090 111.840 ;
        RECT 4.400 105.040 430.090 106.440 ;
        RECT 3.990 96.240 430.090 105.040 ;
        RECT 3.990 94.840 429.690 96.240 ;
        RECT 3.990 89.440 430.090 94.840 ;
        RECT 4.400 88.040 430.090 89.440 ;
        RECT 3.990 79.240 430.090 88.040 ;
        RECT 3.990 77.840 429.690 79.240 ;
        RECT 3.990 72.440 430.090 77.840 ;
        RECT 4.400 71.040 430.090 72.440 ;
        RECT 3.990 58.840 430.090 71.040 ;
        RECT 3.990 57.440 429.690 58.840 ;
        RECT 3.990 52.040 430.090 57.440 ;
        RECT 4.400 50.640 430.090 52.040 ;
        RECT 3.990 41.840 430.090 50.640 ;
        RECT 3.990 40.440 429.690 41.840 ;
        RECT 3.990 35.040 430.090 40.440 ;
        RECT 4.400 33.640 430.090 35.040 ;
        RECT 3.990 24.840 430.090 33.640 ;
        RECT 3.990 23.440 429.690 24.840 ;
        RECT 3.990 18.040 430.090 23.440 ;
        RECT 4.400 16.640 430.090 18.040 ;
        RECT 3.990 4.440 430.090 16.640 ;
        RECT 3.990 3.575 429.690 4.440 ;
      LAYER met4 ;
        RECT 68.375 11.735 174.240 430.945 ;
        RECT 176.640 11.735 177.540 430.945 ;
        RECT 179.940 11.735 327.840 430.945 ;
        RECT 330.240 11.735 331.140 430.945 ;
        RECT 333.540 11.735 371.385 430.945 ;
  END
END alu_32_bit
END LIBRARY


magic
tech sky130A
magscale 1 2
timestamp 1752826596
<< obsli1 >>
rect 1104 2159 85652 86513
<< obsm1 >>
rect 14 2128 85730 86544
<< metal2 >>
rect 18 88162 74 88962
rect 3238 88162 3294 88962
rect 7102 88162 7158 88962
rect 10322 88162 10378 88962
rect 13542 88162 13598 88962
rect 17406 88162 17462 88962
rect 20626 88162 20682 88962
rect 23846 88162 23902 88962
rect 27066 88162 27122 88962
rect 30930 88162 30986 88962
rect 34150 88162 34206 88962
rect 37370 88162 37426 88962
rect 40590 88162 40646 88962
rect 44454 88162 44510 88962
rect 47674 88162 47730 88962
rect 50894 88162 50950 88962
rect 54114 88162 54170 88962
rect 57978 88162 58034 88962
rect 61198 88162 61254 88962
rect 64418 88162 64474 88962
rect 68282 88162 68338 88962
rect 71502 88162 71558 88962
rect 74722 88162 74778 88962
rect 77942 88162 77998 88962
rect 81806 88162 81862 88962
rect 85026 88162 85082 88962
rect 18 0 74 800
rect 3238 0 3294 800
rect 6458 0 6514 800
rect 9678 0 9734 800
rect 13542 0 13598 800
rect 16762 0 16818 800
rect 19982 0 20038 800
rect 23202 0 23258 800
rect 27066 0 27122 800
rect 30286 0 30342 800
rect 33506 0 33562 800
rect 36726 0 36782 800
rect 40590 0 40646 800
rect 43810 0 43866 800
rect 47030 0 47086 800
rect 50894 0 50950 800
rect 54114 0 54170 800
rect 57334 0 57390 800
rect 60554 0 60610 800
rect 64418 0 64474 800
rect 67638 0 67694 800
rect 70858 0 70914 800
rect 74078 0 74134 800
rect 77942 0 77998 800
rect 81162 0 81218 800
rect 84382 0 84438 800
<< obsm2 >>
rect 130 88106 3182 88162
rect 3350 88106 7046 88162
rect 7214 88106 10266 88162
rect 10434 88106 13486 88162
rect 13654 88106 17350 88162
rect 17518 88106 20570 88162
rect 20738 88106 23790 88162
rect 23958 88106 27010 88162
rect 27178 88106 30874 88162
rect 31042 88106 34094 88162
rect 34262 88106 37314 88162
rect 37482 88106 40534 88162
rect 40702 88106 44398 88162
rect 44566 88106 47618 88162
rect 47786 88106 50838 88162
rect 51006 88106 54058 88162
rect 54226 88106 57922 88162
rect 58090 88106 61142 88162
rect 61310 88106 64362 88162
rect 64530 88106 68226 88162
rect 68394 88106 71446 88162
rect 71614 88106 74666 88162
rect 74834 88106 77886 88162
rect 78054 88106 81750 88162
rect 81918 88106 84970 88162
rect 85138 88106 85726 88162
rect 20 856 85726 88106
rect 130 711 3182 856
rect 3350 711 6402 856
rect 6570 711 9622 856
rect 9790 711 13486 856
rect 13654 711 16706 856
rect 16874 711 19926 856
rect 20094 711 23146 856
rect 23314 711 27010 856
rect 27178 711 30230 856
rect 30398 711 33450 856
rect 33618 711 36670 856
rect 36838 711 40534 856
rect 40702 711 43754 856
rect 43922 711 46974 856
rect 47142 711 50838 856
rect 51006 711 54058 856
rect 54226 711 57278 856
rect 57446 711 60498 856
rect 60666 711 64362 856
rect 64530 711 67582 856
rect 67750 711 70802 856
rect 70970 711 74022 856
rect 74190 711 77886 856
rect 78054 711 81106 856
rect 81274 711 84326 856
rect 84494 711 85726 856
<< metal3 >>
rect 86018 87048 86818 87168
rect 0 85688 800 85808
rect 86018 83648 86818 83768
rect 0 82288 800 82408
rect 86018 79568 86818 79688
rect 0 78208 800 78328
rect 86018 76168 86818 76288
rect 0 74808 800 74928
rect 86018 72768 86818 72888
rect 0 71408 800 71528
rect 86018 69368 86818 69488
rect 0 68008 800 68128
rect 86018 65288 86818 65408
rect 0 63928 800 64048
rect 86018 61888 86818 62008
rect 0 60528 800 60648
rect 86018 58488 86818 58608
rect 0 57128 800 57248
rect 86018 54408 86818 54528
rect 0 53728 800 53848
rect 86018 51008 86818 51128
rect 0 49648 800 49768
rect 86018 47608 86818 47728
rect 0 46248 800 46368
rect 86018 44208 86818 44328
rect 0 42848 800 42968
rect 86018 40128 86818 40248
rect 0 38768 800 38888
rect 86018 36728 86818 36848
rect 0 35368 800 35488
rect 86018 33328 86818 33448
rect 0 31968 800 32088
rect 86018 29928 86818 30048
rect 0 28568 800 28688
rect 86018 25848 86818 25968
rect 0 24488 800 24608
rect 86018 22448 86818 22568
rect 0 21088 800 21208
rect 86018 19048 86818 19168
rect 0 17688 800 17808
rect 86018 15648 86818 15768
rect 0 14288 800 14408
rect 86018 11568 86818 11688
rect 0 10208 800 10328
rect 86018 8168 86818 8288
rect 0 6808 800 6928
rect 86018 4768 86818 4888
rect 0 3408 800 3528
rect 86018 688 86818 808
<< obsm3 >>
rect 798 86968 85938 87141
rect 798 85888 86018 86968
rect 880 85608 86018 85888
rect 798 83848 86018 85608
rect 798 83568 85938 83848
rect 798 82488 86018 83568
rect 880 82208 86018 82488
rect 798 79768 86018 82208
rect 798 79488 85938 79768
rect 798 78408 86018 79488
rect 880 78128 86018 78408
rect 798 76368 86018 78128
rect 798 76088 85938 76368
rect 798 75008 86018 76088
rect 880 74728 86018 75008
rect 798 72968 86018 74728
rect 798 72688 85938 72968
rect 798 71608 86018 72688
rect 880 71328 86018 71608
rect 798 69568 86018 71328
rect 798 69288 85938 69568
rect 798 68208 86018 69288
rect 880 67928 86018 68208
rect 798 65488 86018 67928
rect 798 65208 85938 65488
rect 798 64128 86018 65208
rect 880 63848 86018 64128
rect 798 62088 86018 63848
rect 798 61808 85938 62088
rect 798 60728 86018 61808
rect 880 60448 86018 60728
rect 798 58688 86018 60448
rect 798 58408 85938 58688
rect 798 57328 86018 58408
rect 880 57048 86018 57328
rect 798 54608 86018 57048
rect 798 54328 85938 54608
rect 798 53928 86018 54328
rect 880 53648 86018 53928
rect 798 51208 86018 53648
rect 798 50928 85938 51208
rect 798 49848 86018 50928
rect 880 49568 86018 49848
rect 798 47808 86018 49568
rect 798 47528 85938 47808
rect 798 46448 86018 47528
rect 880 46168 86018 46448
rect 798 44408 86018 46168
rect 798 44128 85938 44408
rect 798 43048 86018 44128
rect 880 42768 86018 43048
rect 798 40328 86018 42768
rect 798 40048 85938 40328
rect 798 38968 86018 40048
rect 880 38688 86018 38968
rect 798 36928 86018 38688
rect 798 36648 85938 36928
rect 798 35568 86018 36648
rect 880 35288 86018 35568
rect 798 33528 86018 35288
rect 798 33248 85938 33528
rect 798 32168 86018 33248
rect 880 31888 86018 32168
rect 798 30128 86018 31888
rect 798 29848 85938 30128
rect 798 28768 86018 29848
rect 880 28488 86018 28768
rect 798 26048 86018 28488
rect 798 25768 85938 26048
rect 798 24688 86018 25768
rect 880 24408 86018 24688
rect 798 22648 86018 24408
rect 798 22368 85938 22648
rect 798 21288 86018 22368
rect 880 21008 86018 21288
rect 798 19248 86018 21008
rect 798 18968 85938 19248
rect 798 17888 86018 18968
rect 880 17608 86018 17888
rect 798 15848 86018 17608
rect 798 15568 85938 15848
rect 798 14488 86018 15568
rect 880 14208 86018 14488
rect 798 11768 86018 14208
rect 798 11488 85938 11768
rect 798 10408 86018 11488
rect 880 10128 86018 10408
rect 798 8368 86018 10128
rect 798 8088 85938 8368
rect 798 7008 86018 8088
rect 880 6728 86018 7008
rect 798 4968 86018 6728
rect 798 4688 85938 4968
rect 798 3608 86018 4688
rect 880 3328 86018 3608
rect 798 888 86018 3328
rect 798 715 85938 888
<< metal4 >>
rect 4208 2128 4528 86544
rect 4868 2128 5188 86544
rect 34928 2128 35248 86544
rect 35588 2128 35908 86544
rect 65648 2128 65968 86544
rect 66308 2128 66628 86544
<< obsm4 >>
rect 13675 2347 34848 86189
rect 35328 2347 35508 86189
rect 35988 2347 65568 86189
rect 66048 2347 66228 86189
rect 66708 2347 74277 86189
<< metal5 >>
rect 1056 67278 85700 67598
rect 1056 66618 85700 66938
rect 1056 36642 85700 36962
rect 1056 35982 85700 36302
rect 1056 6006 85700 6326
rect 1056 5346 85700 5666
<< labels >>
rlabel metal3 s 86018 87048 86818 87168 6 A[0]
port 1 nsew signal input
rlabel metal3 s 86018 83648 86818 83768 6 A[10]
port 2 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 A[11]
port 3 nsew signal input
rlabel metal3 s 0 60528 800 60648 6 A[12]
port 4 nsew signal input
rlabel metal3 s 0 82288 800 82408 6 A[13]
port 5 nsew signal input
rlabel metal3 s 86018 58488 86818 58608 6 A[14]
port 6 nsew signal input
rlabel metal3 s 86018 29928 86818 30048 6 A[15]
port 7 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 A[16]
port 8 nsew signal input
rlabel metal3 s 86018 11568 86818 11688 6 A[17]
port 9 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 A[18]
port 10 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 A[19]
port 11 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 A[1]
port 12 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 A[20]
port 13 nsew signal input
rlabel metal2 s 57978 88162 58034 88962 6 A[21]
port 14 nsew signal input
rlabel metal2 s 20626 88162 20682 88962 6 A[22]
port 15 nsew signal input
rlabel metal2 s 23846 88162 23902 88962 6 A[23]
port 16 nsew signal input
rlabel metal3 s 86018 47608 86818 47728 6 A[24]
port 17 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 A[25]
port 18 nsew signal input
rlabel metal3 s 86018 79568 86818 79688 6 A[26]
port 19 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 A[27]
port 20 nsew signal input
rlabel metal3 s 86018 65288 86818 65408 6 A[28]
port 21 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 A[29]
port 22 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 A[2]
port 23 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 A[30]
port 24 nsew signal input
rlabel metal2 s 54114 88162 54170 88962 6 A[31]
port 25 nsew signal input
rlabel metal3 s 86018 44208 86818 44328 6 A[3]
port 26 nsew signal input
rlabel metal2 s 30930 88162 30986 88962 6 A[4]
port 27 nsew signal input
rlabel metal2 s 34150 88162 34206 88962 6 A[5]
port 28 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 A[6]
port 29 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 A[7]
port 30 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 A[8]
port 31 nsew signal input
rlabel metal3 s 86018 76168 86818 76288 6 A[9]
port 32 nsew signal input
rlabel metal3 s 86018 19048 86818 19168 6 B[0]
port 33 nsew signal input
rlabel metal2 s 50894 88162 50950 88962 6 B[10]
port 34 nsew signal input
rlabel metal3 s 86018 25848 86818 25968 6 B[11]
port 35 nsew signal input
rlabel metal2 s 37370 88162 37426 88962 6 B[12]
port 36 nsew signal input
rlabel metal2 s 64418 88162 64474 88962 6 B[13]
port 37 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 B[14]
port 38 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 B[15]
port 39 nsew signal input
rlabel metal3 s 86018 4768 86818 4888 6 B[16]
port 40 nsew signal input
rlabel metal3 s 86018 72768 86818 72888 6 B[17]
port 41 nsew signal input
rlabel metal3 s 86018 36728 86818 36848 6 B[18]
port 42 nsew signal input
rlabel metal2 s 44454 88162 44510 88962 6 B[19]
port 43 nsew signal input
rlabel metal2 s 71502 88162 71558 88962 6 B[1]
port 44 nsew signal input
rlabel metal3 s 86018 688 86818 808 6 B[20]
port 45 nsew signal input
rlabel metal3 s 86018 69368 86818 69488 6 B[21]
port 46 nsew signal input
rlabel metal2 s 81806 88162 81862 88962 6 B[22]
port 47 nsew signal input
rlabel metal2 s 47674 88162 47730 88962 6 B[23]
port 48 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 B[24]
port 49 nsew signal input
rlabel metal3 s 86018 15648 86818 15768 6 B[25]
port 50 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 B[26]
port 51 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 B[27]
port 52 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 B[28]
port 53 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 B[29]
port 54 nsew signal input
rlabel metal2 s 27066 88162 27122 88962 6 B[2]
port 55 nsew signal input
rlabel metal2 s 74722 88162 74778 88962 6 B[30]
port 56 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 B[31]
port 57 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 B[3]
port 58 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 B[4]
port 59 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 B[5]
port 60 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 B[6]
port 61 nsew signal input
rlabel metal3 s 86018 22448 86818 22568 6 B[7]
port 62 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 B[8]
port 63 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 B[9]
port 64 nsew signal input
rlabel metal4 s 4868 2128 5188 86544 6 VGND
port 65 nsew ground bidirectional
rlabel metal4 s 35588 2128 35908 86544 6 VGND
port 65 nsew ground bidirectional
rlabel metal4 s 66308 2128 66628 86544 6 VGND
port 65 nsew ground bidirectional
rlabel metal5 s 1056 6006 85700 6326 6 VGND
port 65 nsew ground bidirectional
rlabel metal5 s 1056 36642 85700 36962 6 VGND
port 65 nsew ground bidirectional
rlabel metal5 s 1056 67278 85700 67598 6 VGND
port 65 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 86544 6 VPWR
port 66 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 86544 6 VPWR
port 66 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 86544 6 VPWR
port 66 nsew power bidirectional
rlabel metal5 s 1056 5346 85700 5666 6 VPWR
port 66 nsew power bidirectional
rlabel metal5 s 1056 35982 85700 36302 6 VPWR
port 66 nsew power bidirectional
rlabel metal5 s 1056 66618 85700 66938 6 VPWR
port 66 nsew power bidirectional
rlabel metal3 s 0 57128 800 57248 6 control[0]
port 67 nsew signal input
rlabel metal2 s 10322 88162 10378 88962 6 control[1]
port 68 nsew signal input
rlabel metal3 s 86018 33328 86818 33448 6 control[2]
port 69 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 control[3]
port 70 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 result[0]
port 71 nsew signal output
rlabel metal3 s 86018 61888 86818 62008 6 result[10]
port 72 nsew signal output
rlabel metal2 s 13542 88162 13598 88962 6 result[11]
port 73 nsew signal output
rlabel metal3 s 0 53728 800 53848 6 result[12]
port 74 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 result[13]
port 75 nsew signal output
rlabel metal2 s 18 0 74 800 6 result[14]
port 76 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 result[15]
port 77 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 result[16]
port 78 nsew signal output
rlabel metal2 s 40590 88162 40646 88962 6 result[17]
port 79 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 result[18]
port 80 nsew signal output
rlabel metal2 s 18 88162 74 88962 6 result[19]
port 81 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 result[1]
port 82 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 result[20]
port 83 nsew signal output
rlabel metal2 s 77942 88162 77998 88962 6 result[21]
port 84 nsew signal output
rlabel metal2 s 61198 88162 61254 88962 6 result[22]
port 85 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 result[23]
port 86 nsew signal output
rlabel metal2 s 85026 88162 85082 88962 6 result[24]
port 87 nsew signal output
rlabel metal3 s 86018 8168 86818 8288 6 result[25]
port 88 nsew signal output
rlabel metal2 s 3238 88162 3294 88962 6 result[26]
port 89 nsew signal output
rlabel metal3 s 86018 51008 86818 51128 6 result[27]
port 90 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 result[28]
port 91 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 result[29]
port 92 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 result[2]
port 93 nsew signal output
rlabel metal3 s 86018 54408 86818 54528 6 result[30]
port 94 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 result[31]
port 95 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 result[3]
port 96 nsew signal output
rlabel metal2 s 68282 88162 68338 88962 6 result[4]
port 97 nsew signal output
rlabel metal2 s 7102 88162 7158 88962 6 result[5]
port 98 nsew signal output
rlabel metal2 s 17406 88162 17462 88962 6 result[6]
port 99 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 result[7]
port 100 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 result[8]
port 101 nsew signal output
rlabel metal3 s 0 78208 800 78328 6 result[9]
port 102 nsew signal output
rlabel metal3 s 86018 40128 86818 40248 6 zero_flag
port 103 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 86818 88962
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 13072464
string GDS_FILE /openlane/designs/ALU/runs/RUN_2025.07.18_08.04.31/results/signoff/alu_32_bit.magic.gds
string GDS_START 1216130
<< end >>


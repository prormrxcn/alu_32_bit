* NGSPICE file created from alu_32_bit.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

.subckt alu_32_bit A[0] A[10] A[11] A[12] A[13] A[14] A[15] A[16] A[17] A[18] A[19]
+ A[1] A[20] A[21] A[22] A[23] A[24] A[25] A[26] A[27] A[28] A[29] A[2] A[30] A[31]
+ A[3] A[4] A[5] A[6] A[7] A[8] A[9] B[0] B[10] B[11] B[12] B[13] B[14] B[15] B[16]
+ B[17] B[18] B[19] B[1] B[20] B[21] B[22] B[23] B[24] B[25] B[26] B[27] B[28] B[29]
+ B[2] B[30] B[31] B[3] B[4] B[5] B[6] B[7] B[8] B[9] VGND VPWR control[0] control[1]
+ control[2] control[3] result[0] result[10] result[11] result[12] result[13] result[14]
+ result[15] result[16] result[17] result[18] result[19] result[1] result[20] result[21]
+ result[22] result[23] result[24] result[25] result[26] result[27] result[28] result[29]
+ result[2] result[30] result[31] result[3] result[4] result[5] result[6] result[7]
+ result[8] result[9] zero_flag
XFILLER_0_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6914_ net129 _1620_ _1623_ _2492_ VGND VGND VPWR VPWR _2493_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_134_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6845_ _2406_ _2415_ VGND VGND VPWR VPWR _2417_ sky130_fd_sc_hd__nand2_1
X_6776_ _2134_ _2135_ _2133_ VGND VGND VPWR VPWR _2341_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_91_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3988_ _2292_ _2478_ _2631_ _2806_ _0554_ _0183_ VGND VGND VPWR VPWR _2817_ sky130_fd_sc_hd__mux4_1
XFILLER_0_64_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5727_ _1077_ _1084_ VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__or2_2
XFILLER_0_73_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5658_ _1116_ _1117_ _1118_ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__and3_4
XFILLER_0_130_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4609_ _3711_ VGND VGND VPWR VPWR _3712_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5589_ _1041_ _1042_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7328_ _3273_ _1756_ VGND VGND VPWR VPWR _2944_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7259_ _3213_ _0305_ _1309_ _2869_ _0867_ _0573_ VGND VGND VPWR VPWR _2870_ sky130_fd_sc_hd__mux4_1
XFILLER_0_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer7 _3529_ VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__buf_1
XFILLER_0_23_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4960_ _0332_ _0333_ _0354_ _0355_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4891_ _0279_ _0280_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__xnor2_2
X_3911_ _1942_ _1963_ _0892_ VGND VGND VPWR VPWR _1974_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3842_ _1144_ _1154_ _1165_ net65 VGND VGND VPWR VPWR _1220_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_74_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6630_ _3425_ _3513_ _2510_ _2543_ _2039_ VGND VGND VPWR VPWR _2181_ sky130_fd_sc_hd__a41o_1
XFILLER_0_7_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6561_ _1789_ _1786_ _1925_ VGND VGND VPWR VPWR _2107_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3773_ net1 VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__clkbuf_4
X_5512_ _0373_ net7 net8 _3352_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6492_ _1872_ _1880_ VGND VGND VPWR VPWR _2031_ sky130_fd_sc_hd__and2_1
X_5443_ _0883_ _3698_ _0870_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5374_ _0741_ _0742_ _0806_ _0807_ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__a22o_1
X_7113_ _0881_ _0521_ net22 _2051_ VGND VGND VPWR VPWR _2710_ sky130_fd_sc_hd__nand4_2
X_4325_ _3343_ VGND VGND VPWR VPWR _3430_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4256_ _3316_ _3318_ _3317_ VGND VGND VPWR VPWR _3362_ sky130_fd_sc_hd__a21bo_1
X_7044_ _2633_ _2634_ VGND VGND VPWR VPWR _2635_ sky130_fd_sc_hd__or2_1
X_4187_ _3108_ _3293_ VGND VGND VPWR VPWR _3294_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6828_ _2395_ _2396_ _2333_ _2189_ VGND VGND VPWR VPWR _2398_ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6759_ _3730_ _2319_ _2321_ _0575_ VGND VGND VPWR VPWR _2322_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_61_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5090_ _0495_ _0496_ _0492_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__o21ai_1
X_4110_ _0838_ _3126_ _3213_ _3217_ _2980_ VGND VGND VPWR VPWR _3218_ sky130_fd_sc_hd__a32o_1
XFILLER_0_75_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4041_ _1952_ _1745_ _0892_ VGND VGND VPWR VPWR _3150_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5992_ _0335_ net46 net47 _0434_ VGND VGND VPWR VPWR _1484_ sky130_fd_sc_hd__a22o_1
X_4943_ _0205_ _3718_ _0099_ _0335_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_47_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4874_ _0253_ _0261_ _0262_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__nand3_1
XFILLER_0_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6613_ _2151_ _2152_ _2162_ VGND VGND VPWR VPWR _2163_ sky130_fd_sc_hd__or3_4
XFILLER_0_144_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3825_ _0226_ VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__buf_4
XFILLER_0_43_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3756_ net55 VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__buf_8
XFILLER_0_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6544_ _2085_ _2086_ _1903_ _1905_ VGND VGND VPWR VPWR _2088_ sky130_fd_sc_hd__a211o_1
X_6475_ _2006_ _2008_ _2009_ VGND VGND VPWR VPWR _2012_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_43_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5426_ _0862_ _2587_ _3128_ _0558_ _0863_ _0864_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__mux4_1
XFILLER_0_113_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5357_ _0629_ _0631_ _0632_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_100_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4308_ _1187_ VGND VGND VPWR VPWR _3414_ sky130_fd_sc_hd__clkbuf_4
X_5288_ _0573_ _3587_ _0703_ _0709_ _0714_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__a311o_1
X_4239_ net23 net12 net61 net62 VGND VGND VPWR VPWR _3345_ sky130_fd_sc_hd__and4_1
X_7027_ _2615_ VGND VGND VPWR VPWR _2616_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_640 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap5 _1737_ VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_88_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4590_ _3692_ VGND VGND VPWR VPWR _3693_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6260_ _1272_ _1273_ _1300_ VGND VGND VPWR VPWR _1777_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5211_ _3452_ _2489_ _2521_ _3449_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__a22o_1
X_6191_ _0488_ _0390_ net16 net17 VGND VGND VPWR VPWR _1702_ sky130_fd_sc_hd__nand4_2
X_5142_ _0546_ _0555_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5073_ _0476_ _0478_ _0479_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__nand3_4
X_4024_ _2718_ VGND VGND VPWR VPWR _3133_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5975_ _1450_ _1462_ _1463_ _3161_ _1464_ VGND VGND VPWR VPWR _1465_ sky130_fd_sc_hd__a221o_1
X_4926_ _0290_ _0291_ _0319_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__o21ai_4
XFILLER_0_75_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4857_ _0240_ _0243_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__xor2_2
XFILLER_0_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3808_ net66 net68 net67 net65 VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4788_ _0090_ _0076_ _0166_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6527_ _2067_ _2068_ VGND VGND VPWR VPWR _2069_ sky130_fd_sc_hd__xor2_2
XFILLER_0_113_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3739_ _0085_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__buf_4
XFILLER_0_70_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6458_ _0401_ _1767_ net19 _0499_ VGND VGND VPWR VPWR _1993_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5409_ _0428_ _0846_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__or2_1
X_6389_ _1790_ _1746_ _1916_ _1917_ VGND VGND VPWR VPWR _1918_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_98_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire111 _1068_ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__buf_1
XFILLER_0_124_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5760_ _0042_ _2499_ VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__nand2_1
X_4711_ _0081_ _0083_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__and2_1
X_5691_ _1153_ _0995_ _1140_ VGND VGND VPWR VPWR _1155_ sky130_fd_sc_hd__or3_4
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7430_ _0455_ _0696_ VGND VGND VPWR VPWR _3055_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4642_ _3685_ _3137_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__and2b_1
XFILLER_0_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4573_ _3612_ _3674_ _3675_ VGND VGND VPWR VPWR _3676_ sky130_fd_sc_hd__and3_1
XFILLER_0_112_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7361_ _2976_ _2979_ VGND VGND VPWR VPWR _2981_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7292_ _2767_ _2798_ _2904_ VGND VGND VPWR VPWR _2905_ sky130_fd_sc_hd__a21o_1
X_6312_ _1831_ _1833_ _2117_ _0654_ VGND VGND VPWR VPWR _1834_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_12_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6243_ _0004_ _0585_ _1017_ _1758_ _0429_ _0189_ VGND VGND VPWR VPWR _1759_ sky130_fd_sc_hd__mux4_1
XFILLER_0_12_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6174_ _2248_ _2653_ _0339_ _0099_ VGND VGND VPWR VPWR _1683_ sky130_fd_sc_hd__nand4_4
X_5125_ _0533_ _0534_ _0535_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5056_ _0450_ _0460_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4007_ _0554_ _0936_ VGND VGND VPWR VPWR _3024_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5958_ _1295_ _1942_ VGND VGND VPWR VPWR _1446_ sky130_fd_sc_hd__and2b_1
XFILLER_0_75_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4909_ _0175_ _0186_ _0296_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5889_ _3511_ _0491_ _2686_ _0104_ VGND VGND VPWR VPWR _1371_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_5 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer17 net140 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6930_ _2337_ _2338_ _2336_ VGND VGND VPWR VPWR _2509_ sky130_fd_sc_hd__a21bo_1
Xrebuffer28 _2147_ VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_1
Xrebuffer39 net204 VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__buf_2
XFILLER_0_88_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6861_ _2431_ _2432_ _2418_ VGND VGND VPWR VPWR _2435_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6792_ _3272_ _1898_ _1931_ _3197_ VGND VGND VPWR VPWR _2359_ sky130_fd_sc_hd__a22o_1
X_5812_ _3155_ _1287_ _0861_ VGND VGND VPWR VPWR _1288_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5743_ _1202_ _1211_ VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__xor2_1
XFILLER_0_18_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5674_ _0897_ _0989_ _0988_ VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_5_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4625_ _3580_ VGND VGND VPWR VPWR _3727_ sky130_fd_sc_hd__buf_2
XFILLER_0_5_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7413_ _2857_ _3037_ VGND VGND VPWR VPWR _3038_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4556_ _3649_ _3657_ _3658_ VGND VGND VPWR VPWR _3659_ sky130_fd_sc_hd__nand3_1
XFILLER_0_115_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7344_ _3135_ _0559_ VGND VGND VPWR VPWR _2962_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4487_ _0969_ VGND VGND VPWR VPWR _3591_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7275_ _2884_ _2885_ VGND VGND VPWR VPWR _2886_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6226_ net108 _1738_ _1577_ _1579_ VGND VGND VPWR VPWR _1740_ sky130_fd_sc_hd__o211a_4
X_6157_ _2445_ _0688_ _1662_ _1663_ VGND VGND VPWR VPWR _1664_ sky130_fd_sc_hd__nand4_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _0377_ _0387_ _0386_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__a21bo_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6088_ _1586_ _1587_ _1480_ VGND VGND VPWR VPWR _1589_ sky130_fd_sc_hd__a21o_1
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5039_ _3571_ _0427_ _0432_ _0442_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__a211o_1
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput75 net75 VGND VGND VPWR VPWR result[15] sky130_fd_sc_hd__clkbuf_4
Xoutput97 net97 VGND VGND VPWR VPWR result[6] sky130_fd_sc_hd__clkbuf_4
Xoutput86 net86 VGND VGND VPWR VPWR result[25] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4410_ _0445_ _3424_ _3513_ _0991_ VGND VGND VPWR VPWR _3514_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_2_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5390_ _2587_ _0722_ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__and2_2
XFILLER_0_111_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4341_ _3441_ _3445_ VGND VGND VPWR VPWR _3446_ sky130_fd_sc_hd__xor2_2
XFILLER_0_50_782 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4272_ net186 _3375_ net196 VGND VGND VPWR VPWR _3378_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_10_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7060_ _2610_ _2611_ _2649_ _2650_ VGND VGND VPWR VPWR _2652_ sky130_fd_sc_hd__a22o_1
X_6011_ _2390_ _0688_ _1502_ _1503_ VGND VGND VPWR VPWR _1505_ sky130_fd_sc_hd__nand4_1
XFILLER_0_118_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6913_ _1754_ _1926_ _2105_ _2275_ VGND VGND VPWR VPWR _2492_ sky130_fd_sc_hd__or4_4
XFILLER_0_49_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6844_ _2406_ _2415_ VGND VGND VPWR VPWR _2416_ sky130_fd_sc_hd__or2_2
X_6775_ _2336_ _2337_ _2338_ VGND VGND VPWR VPWR _2340_ sky130_fd_sc_hd__a21o_1
X_3987_ _2729_ _2795_ _0936_ VGND VGND VPWR VPWR _2806_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5726_ _1083_ _1082_ VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__or2b_1
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_532 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5657_ _0962_ _0971_ _0970_ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_5_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4608_ _1165_ _0630_ _1144_ _1154_ VGND VGND VPWR VPWR _3711_ sky130_fd_sc_hd__or4b_1
X_5588_ _0466_ _1007_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4539_ _3629_ _3641_ VGND VGND VPWR VPWR _3642_ sky130_fd_sc_hd__xor2_2
X_7327_ _2939_ _2942_ VGND VGND VPWR VPWR _2943_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7258_ _2114_ _2868_ _0866_ VGND VGND VPWR VPWR _2869_ sky130_fd_sc_hd__mux2_1
X_6209_ _1716_ _1717_ _1718_ VGND VGND VPWR VPWR _1721_ sky130_fd_sc_hd__a21oi_2
X_7189_ _2786_ _2792_ VGND VGND VPWR VPWR _2793_ sky130_fd_sc_hd__xnor2_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer8 _0993_ VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4890_ _0092_ _0158_ _0157_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_86_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3910_ _1952_ VGND VGND VPWR VPWR _1963_ sky130_fd_sc_hd__buf_4
XFILLER_0_58_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3841_ _1198_ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__buf_2
XFILLER_0_117_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3772_ _0401_ _0445_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_55_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6560_ _1964_ _2104_ VGND VGND VPWR VPWR _2105_ sky130_fd_sc_hd__xnor2_4
X_5511_ _3352_ _0373_ net7 VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6491_ _1879_ _1873_ VGND VGND VPWR VPWR _2030_ sky130_fd_sc_hd__and2b_1
XFILLER_0_152_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5442_ _0882_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5373_ _0741_ _0742_ _0806_ _0807_ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__nand4_2
XFILLER_0_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4324_ _0205_ _2892_ _3354_ _3353_ _0172_ VGND VGND VPWR VPWR _3429_ sky130_fd_sc_hd__a32o_1
X_7112_ _0521_ net22 net24 _0881_ VGND VGND VPWR VPWR _2709_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7043_ _0226_ _1949_ _2630_ _2632_ VGND VGND VPWR VPWR _2634_ sky130_fd_sc_hd__and4_1
X_4255_ _3358_ _3359_ _3357_ VGND VGND VPWR VPWR _3361_ sky130_fd_sc_hd__a21o_1
X_4186_ _3291_ _3292_ _1712_ VGND VGND VPWR VPWR _3293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6827_ _2333_ _2189_ _2395_ _2396_ VGND VGND VPWR VPWR _2397_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6758_ _0573_ _2073_ _3729_ _2320_ VGND VGND VPWR VPWR _2321_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5709_ _1051_ _1053_ VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__or2_1
X_6689_ _0205_ net49 net50 _0335_ VGND VGND VPWR VPWR _2246_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_590 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_468 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4040_ _1909_ _1942_ _0892_ VGND VGND VPWR VPWR _3149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5991_ _0346_ _0707_ net46 _1294_ VGND VGND VPWR VPWR _1483_ sky130_fd_sc_hd__and4_1
XFILLER_0_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4942_ net38 VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4873_ _0257_ _0258_ _0260_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__a21o_1
X_6612_ _2153_ _2161_ VGND VGND VPWR VPWR _2162_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_144_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3824_ _0117_ VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__buf_4
XFILLER_0_104_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3755_ net55 net23 VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6543_ _1903_ _1905_ _2085_ _2086_ VGND VGND VPWR VPWR _2087_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_43_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6474_ _2010_ VGND VGND VPWR VPWR _2011_ sky130_fd_sc_hd__buf_2
XFILLER_0_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5425_ _0584_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5356_ _0786_ _0787_ _0785_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4307_ _3387_ _3412_ VGND VGND VPWR VPWR _3413_ sky130_fd_sc_hd__nor2_1
X_5287_ _3727_ _0711_ _0713_ _0849_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__o211a_1
X_4238_ net23 net61 _3270_ _0412_ VGND VGND VPWR VPWR _3344_ sky130_fd_sc_hd__a22oi_1
X_7026_ _1045_ net52 _2299_ _1056_ VGND VGND VPWR VPWR _2615_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4169_ _3274_ _3275_ VGND VGND VPWR VPWR _3276_ sky130_fd_sc_hd__or2_2
XFILLER_0_97_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_700 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap6 _0398_ VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5210_ _0292_ _0380_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6190_ _1554_ _1573_ _1574_ VGND VGND VPWR VPWR _1700_ sky130_fd_sc_hd__nor3_1
X_5141_ _0549_ _0552_ _0553_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__and3_1
X_5072_ _0095_ _0110_ _0348_ _0347_ _3423_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__a32o_1
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4023_ _3129_ _3130_ _3131_ VGND VGND VPWR VPWR _3132_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5974_ _3712_ _1450_ _1451_ _0309_ VGND VGND VPWR VPWR _1464_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_136_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_755 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4925_ _0181_ _0299_ _0300_ _0318_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__o31a_2
XFILLER_0_59_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4856_ _3632_ _0241_ _0242_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3807_ _0827_ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__buf_4
XFILLER_0_62_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4787_ _0167_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6526_ _1822_ _1824_ VGND VGND VPWR VPWR _2068_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3738_ _0074_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__buf_2
XFILLER_0_43_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6457_ _0499_ _0401_ _1767_ _1799_ VGND VGND VPWR VPWR _1992_ sky130_fd_sc_hd__nand4_1
X_5408_ _3207_ _3602_ _0304_ _0845_ _0429_ _0189_ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__mux4_1
X_6388_ _1914_ _1915_ _1813_ VGND VGND VPWR VPWR _1917_ sky130_fd_sc_hd__a21o_1
X_5339_ _0624_ _0625_ _0626_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_98_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7009_ _2594_ _2595_ VGND VGND VPWR VPWR _2596_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4710_ _0081_ net142 VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__nor2_1
X_5690_ _0814_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4641_ _3721_ _0001_ _0009_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_142_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4572_ _3672_ _3673_ net144 _3611_ VGND VGND VPWR VPWR _3675_ sky130_fd_sc_hd__o211ai_4
X_7360_ _2977_ _2978_ VGND VGND VPWR VPWR _2979_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7291_ _2768_ _2797_ VGND VGND VPWR VPWR _2904_ sky130_fd_sc_hd__nor2_1
X_6311_ _2204_ _0326_ _0453_ _0247_ VGND VGND VPWR VPWR _1833_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6242_ _1756_ _1963_ _1942_ _1909_ _0583_ _0584_ VGND VGND VPWR VPWR _1758_ sky130_fd_sc_hd__mux4_1
XFILLER_0_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6173_ _0491_ _0339_ _0099_ _2248_ VGND VGND VPWR VPWR _1682_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5124_ _0533_ _0534_ _0535_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5055_ _0458_ _0459_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__nor2_1
X_4006_ _2936_ _2991_ VGND VGND VPWR VPWR _3013_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5957_ _3571_ _1302_ _1303_ _1316_ _1445_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__a311o_4
XFILLER_0_137_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4908_ _0296_ _0298_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5888_ _3423_ _0105_ _0491_ _2696_ VGND VGND VPWR VPWR _1370_ sky130_fd_sc_hd__nand4_1
XFILLER_0_63_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4839_ _0085_ _2302_ _3422_ _3572_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__and4_1
XFILLER_0_51_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7489_ net70 net71 _3115_ VGND VGND VPWR VPWR _3116_ sky130_fd_sc_hd__or3_1
X_6509_ _2027_ _2028_ _2047_ _2048_ VGND VGND VPWR VPWR _2049_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_30_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_438 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_6 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer18 _0083_ VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer29 _1619_ VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6860_ _2418_ _2431_ _2432_ VGND VGND VPWR VPWR _2433_ sky130_fd_sc_hd__nand3_2
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6791_ _3197_ _3273_ _1898_ _1931_ VGND VGND VPWR VPWR _2358_ sky130_fd_sc_hd__nand4_2
X_5811_ _0844_ _1285_ VGND VGND VPWR VPWR _1287_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5742_ _1207_ _1210_ VGND VGND VPWR VPWR _1211_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5673_ _1132_ net161 _1033_ _1035_ VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4624_ _3687_ _3696_ _3723_ _3725_ VGND VGND VPWR VPWR _3726_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_53_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7412_ _3034_ _3036_ VGND VGND VPWR VPWR _3037_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4555_ _3654_ _3655_ _3656_ VGND VGND VPWR VPWR _3658_ sky130_fd_sc_hd__a21o_1
X_7343_ _2819_ _2960_ VGND VGND VPWR VPWR _2961_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4486_ _3589_ _3573_ _3204_ VGND VGND VPWR VPWR _3590_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_12_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7274_ _2871_ _2700_ _2883_ _3596_ VGND VGND VPWR VPWR _2885_ sky130_fd_sc_hd__a31o_1
X_6225_ _1577_ _1579_ net108 _1738_ VGND VGND VPWR VPWR _1739_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6156_ _0247_ _0326_ _0453_ _2117_ VGND VGND VPWR VPWR _1663_ sky130_fd_sc_hd__a22o_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _0514_ _0515_ _0506_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6087_ _1480_ _1586_ _1587_ VGND VGND VPWR VPWR _1588_ sky130_fd_sc_hd__nand3_2
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5038_ _0007_ _0436_ _0437_ _0441_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__a211o_1
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6989_ _2572_ net48 _2401_ _2570_ VGND VGND VPWR VPWR _2574_ sky130_fd_sc_hd__and4b_1
XFILLER_0_91_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput76 net76 VGND VGND VPWR VPWR result[16] sky130_fd_sc_hd__clkbuf_4
Xoutput87 net166 VGND VGND VPWR VPWR result[26] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput98 net98 VGND VGND VPWR VPWR result[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4340_ _3442_ _3443_ _3444_ VGND VGND VPWR VPWR _3445_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_50_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4271_ _3374_ _3375_ _3376_ VGND VGND VPWR VPWR _3377_ sky130_fd_sc_hd__and3_4
XFILLER_0_10_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6010_ _3644_ _0326_ _0453_ _3530_ VGND VGND VPWR VPWR _1503_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6912_ _2326_ _2490_ VGND VGND VPWR VPWR _2491_ sky130_fd_sc_hd__xor2_1
XFILLER_0_134_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_636 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6843_ _2413_ _2414_ VGND VGND VPWR VPWR _2415_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6774_ _2336_ _2337_ _2338_ VGND VGND VPWR VPWR _2339_ sky130_fd_sc_hd__nand3_1
XFILLER_0_92_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3986_ _2762_ _2784_ _2029_ VGND VGND VPWR VPWR _2795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5725_ _1189_ _1190_ _1159_ VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5656_ _1114_ _1115_ _1106_ VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4607_ net124 _3687_ _3204_ VGND VGND VPWR VPWR _3710_ sky130_fd_sc_hd__a21o_1
XFILLER_0_130_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5587_ _1039_ _1040_ VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4538_ _3639_ _3640_ VGND VGND VPWR VPWR _3641_ sky130_fd_sc_hd__nor2_2
X_7326_ _2940_ _2941_ VGND VGND VPWR VPWR _2942_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4469_ net2 _3572_ VGND VGND VPWR VPWR _3573_ sky130_fd_sc_hd__and2_4
X_7257_ _2051_ _2018_ _2007_ _1821_ _0863_ _0864_ VGND VGND VPWR VPWR _2868_ sky130_fd_sc_hd__mux4_1
X_6208_ _1719_ VGND VGND VPWR VPWR _1720_ sky130_fd_sc_hd__clkbuf_2
X_7188_ _2787_ _2791_ VGND VGND VPWR VPWR _2792_ sky130_fd_sc_hd__xor2_1
XFILLER_0_99_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6139_ _1498_ _1511_ _1512_ VGND VGND VPWR VPWR _1644_ sky130_fd_sc_hd__and3_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer9 net132 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3840_ net66 net65 net68 net67 VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__or4b_1
XFILLER_0_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3771_ _0434_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__buf_4
XFILLER_0_39_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5510_ _2881_ _2751_ VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6490_ _1893_ _1901_ VGND VGND VPWR VPWR _2028_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5441_ _3296_ _3292_ _0980_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5372_ net112 _0804_ _0743_ _0744_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_23_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4323_ _3345_ _3347_ VGND VGND VPWR VPWR _3428_ sky130_fd_sc_hd__or2_2
X_7111_ _2522_ _2523_ _2533_ VGND VGND VPWR VPWR _2708_ sky130_fd_sc_hd__nor3_2
XFILLER_0_10_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7042_ _0226_ _1949_ _2630_ _2632_ VGND VGND VPWR VPWR _2633_ sky130_fd_sc_hd__a22oi_1
X_4254_ _3357_ _3358_ _3359_ VGND VGND VPWR VPWR _3360_ sky130_fd_sc_hd__nand3_1
X_4185_ _3150_ _3146_ _0521_ VGND VGND VPWR VPWR _3292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6826_ _2369_ _2370_ _2393_ _2394_ VGND VGND VPWR VPWR _2396_ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_0_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6757_ _0199_ _0428_ _3163_ _0571_ VGND VGND VPWR VPWR _2320_ sky130_fd_sc_hd__o31a_1
XFILLER_0_18_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3969_ _2598_ VGND VGND VPWR VPWR _2609_ sky130_fd_sc_hd__buf_4
X_5708_ _1049_ _1057_ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6688_ _2057_ _2059_ VGND VGND VPWR VPWR _2245_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5639_ _1096_ _1097_ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7309_ _2744_ _2747_ _2745_ VGND VGND VPWR VPWR _2923_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_13_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5990_ _1338_ _1350_ _1352_ VGND VGND VPWR VPWR _1481_ sky130_fd_sc_hd__nor3_2
X_4941_ _0238_ _0245_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4872_ _0257_ _0258_ _0260_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__nand3_1
XFILLER_0_47_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3823_ _0980_ _1002_ VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__nand2_2
X_6611_ _2154_ _2159_ VGND VGND VPWR VPWR _2161_ sky130_fd_sc_hd__xor2_2
XFILLER_0_117_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3754_ _0237_ _0248_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6542_ _2082_ _2083_ _2070_ VGND VGND VPWR VPWR _2086_ sky130_fd_sc_hd__a21o_1
X_6473_ _2006_ _2008_ _2009_ VGND VGND VPWR VPWR _2010_ sky130_fd_sc_hd__and3_1
XFILLER_0_112_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5424_ _0583_ VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__buf_4
XFILLER_0_113_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5355_ _0785_ _0786_ _0787_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__nand3_1
XFILLER_0_57_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4306_ _1209_ _3388_ _3204_ VGND VGND VPWR VPWR _3412_ sky130_fd_sc_hd__o21ba_1
X_5286_ _3727_ _0712_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4237_ net63 VGND VGND VPWR VPWR _3343_ sky130_fd_sc_hd__buf_2
X_7025_ _2449_ VGND VGND VPWR VPWR _2614_ sky130_fd_sc_hd__inv_2
X_4168_ _2456_ _3273_ VGND VGND VPWR VPWR _3275_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4099_ _2412_ _2346_ _1023_ _1034_ _0925_ _3131_ VGND VGND VPWR VPWR _3207_ sky130_fd_sc_hd__mux4_2
XFILLER_0_78_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6809_ _2375_ _0293_ _2762_ _2376_ VGND VGND VPWR VPWR _2377_ sky130_fd_sc_hd__and4b_1
XFILLER_0_37_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_439 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap7 _1420_ VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_639 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5140_ _0288_ _0551_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5071_ _2324_ _0110_ _0474_ _0475_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__a22o_1
X_4022_ _0947_ VGND VGND VPWR VPWR _3131_ sky130_fd_sc_hd__buf_4
XFILLER_0_126_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5973_ _3490_ _0863_ _0864_ _0199_ VGND VGND VPWR VPWR _1463_ sky130_fd_sc_hd__o31a_1
XFILLER_0_149_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4924_ _0301_ _0302_ _0317_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4855_ _2423_ net162 net31 _3433_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4786_ _0090_ _0076_ _0166_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__or3_1
X_3806_ _0052_ VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_439 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3737_ net27 VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__buf_8
XFILLER_0_55_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6525_ _2065_ _2066_ VGND VGND VPWR VPWR _2067_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_42_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6456_ _1870_ _1871_ _1881_ VGND VGND VPWR VPWR _1991_ sky130_fd_sc_hd__nor3_1
XFILLER_0_113_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5407_ _2587_ _3128_ _0558_ _3135_ _0583_ _0584_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6387_ _1813_ _1914_ net185 VGND VGND VPWR VPWR _1916_ sky130_fd_sc_hd__nand3_2
X_5338_ _0617_ _0618_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__or2_1
X_7008_ _2592_ _2593_ _2375_ _2377_ VGND VGND VPWR VPWR _2595_ sky130_fd_sc_hd__a211o_1
X_5269_ _0559_ _0558_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__and2b_1
XFILLER_0_98_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4640_ _3201_ _0002_ _0006_ _0007_ _0008_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4571_ net144 _3611_ _3672_ _3673_ VGND VGND VPWR VPWR _3674_ sky130_fd_sc_hd__a211o_1
XFILLER_0_107_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6310_ _0247_ _2204_ _0326_ _0453_ VGND VGND VPWR VPWR _1831_ sky130_fd_sc_hd__and4_1
XFILLER_0_24_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_612 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7290_ _3685_ _0862_ _2752_ _2750_ VGND VGND VPWR VPWR _2902_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6241_ _1625_ _1754_ _1755_ VGND VGND VPWR VPWR _1757_ sky130_fd_sc_hd__a21boi_1
X_6172_ _1544_ _1552_ _1551_ VGND VGND VPWR VPWR _1681_ sky130_fd_sc_hd__a21o_1
X_5123_ _0322_ _0330_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__and2_1
X_5054_ _0456_ _0457_ _0451_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__a21oi_1
X_4005_ _2936_ _2991_ VGND VGND VPWR VPWR _3002_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5956_ _0320_ _1443_ _1444_ VGND VGND VPWR VPWR _1445_ sky130_fd_sc_hd__and3_1
XFILLER_0_87_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4907_ _0296_ _0298_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__nor2_1
X_5887_ _1367_ _1368_ VGND VGND VPWR VPWR _1369_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_145_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4838_ _3635_ _0104_ _0105_ _3440_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_75_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4769_ _0145_ _0146_ _0147_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__nand3_2
XFILLER_0_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7488_ net99 net100 _3114_ VGND VGND VPWR VPWR _3115_ sky130_fd_sc_hd__or3_1
XFILLER_0_70_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6508_ _2030_ _2031_ _2046_ VGND VGND VPWR VPWR _2048_ sky130_fd_sc_hd__nor3_2
XFILLER_0_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6439_ _0346_ _1607_ net50 _0707_ VGND VGND VPWR VPWR _1972_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_113_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_7 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer19 _2047_ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__buf_1
XFILLER_0_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6790_ _2892_ _1931_ _2143_ _2142_ _1745_ VGND VGND VPWR VPWR _2356_ sky130_fd_sc_hd__a32o_1
XFILLER_0_76_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5810_ _0188_ _1284_ _0189_ VGND VGND VPWR VPWR _1285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5741_ _2160_ _3620_ _1080_ _1208_ VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__a31o_1
XFILLER_0_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5672_ _1033_ _1035_ _1132_ _1134_ VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7411_ _2412_ _1797_ VGND VGND VPWR VPWR _3036_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4623_ _3596_ _3724_ VGND VGND VPWR VPWR _3725_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4554_ _3654_ _3655_ _3656_ VGND VGND VPWR VPWR _3657_ sky130_fd_sc_hd__nand3_1
XFILLER_0_103_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7342_ _2785_ _2796_ _2959_ VGND VGND VPWR VPWR _2960_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7273_ _2871_ _2700_ _2883_ VGND VGND VPWR VPWR _2884_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4485_ _1209_ VGND VGND VPWR VPWR _3589_ sky130_fd_sc_hd__clkbuf_4
X_6224_ _1698_ _1699_ _1735_ _1736_ VGND VGND VPWR VPWR _1738_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6155_ _2117_ _2160_ _0326_ _0453_ VGND VGND VPWR VPWR _1662_ sky130_fd_sc_hd__nand4_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _0506_ _0514_ _0515_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__nand3_2
XFILLER_0_57_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6086_ _1584_ _1585_ net154 _1424_ VGND VGND VPWR VPWR _1587_ sky130_fd_sc_hd__o211ai_2
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5037_ _0421_ _0440_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__nor2_1
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6988_ _2401_ _1448_ _2571_ _2572_ VGND VGND VPWR VPWR _2573_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_153_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5939_ _1254_ _1324_ _1424_ _1425_ VGND VGND VPWR VPWR _1426_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput77 net77 VGND VGND VPWR VPWR result[17] sky130_fd_sc_hd__clkbuf_4
Xoutput88 net88 VGND VGND VPWR VPWR result[27] sky130_fd_sc_hd__clkbuf_4
Xoutput99 net99 VGND VGND VPWR VPWR result[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_718 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4270_ net193 _3332_ _3331_ VGND VGND VPWR VPWR _3376_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6911_ _2487_ _2488_ VGND VGND VPWR VPWR _2490_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6842_ _2409_ _2410_ _2411_ VGND VGND VPWR VPWR _2414_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6773_ _0303_ _1799_ VGND VGND VPWR VPWR _2338_ sky130_fd_sc_hd__and2_1
X_3985_ _2773_ VGND VGND VPWR VPWR _2784_ sky130_fd_sc_hd__buf_4
XFILLER_0_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5724_ _1159_ _1189_ _1190_ VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__nor3_1
XFILLER_0_17_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5655_ _1106_ _1114_ _1115_ VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__nand3_1
XFILLER_0_73_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4606_ _2248_ net35 VGND VGND VPWR VPWR _3709_ sky130_fd_sc_hd__and2_2
XFILLER_0_5_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7325_ _2714_ _2722_ VGND VGND VPWR VPWR _2941_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_559 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5586_ _0335_ _0434_ _0721_ _0874_ VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__nand4_1
XFILLER_0_130_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4537_ _3637_ _3638_ _3630_ VGND VGND VPWR VPWR _3640_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4468_ net34 VGND VGND VPWR VPWR _3572_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7256_ _2863_ _2865_ _2866_ VGND VGND VPWR VPWR _2867_ sky130_fd_sc_hd__a21oi_1
X_6207_ _1716_ _1717_ _1718_ VGND VGND VPWR VPWR _1719_ sky130_fd_sc_hd__and3_1
X_7187_ _2789_ _2790_ VGND VGND VPWR VPWR _2791_ sky130_fd_sc_hd__xor2_1
X_4399_ _1209_ _3480_ _3204_ VGND VGND VPWR VPWR _3504_ sky130_fd_sc_hd__o21ba_1
X_6138_ _1511_ VGND VGND VPWR VPWR _1643_ sky130_fd_sc_hd__inv_2
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6069_ _1566_ _1567_ VGND VGND VPWR VPWR _1568_ sky130_fd_sc_hd__xor2_1
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_383 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_751 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3770_ _0423_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__buf_4
XFILLER_0_54_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5440_ _0826_ _0836_ _0878_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__or3b_1
XFILLER_0_15_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5371_ _0743_ _0744_ net112 _0804_ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__a211o_4
XFILLER_0_10_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4322_ _3421_ _3426_ VGND VGND VPWR VPWR _3427_ sky130_fd_sc_hd__xnor2_2
X_7110_ _2536_ _2537_ _2560_ _2561_ VGND VGND VPWR VPWR _2706_ sky130_fd_sc_hd__and4_1
XFILLER_0_10_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4253_ net44 net30 net31 net33 VGND VGND VPWR VPWR _3359_ sky130_fd_sc_hd__a22o_1
X_7041_ _0117_ _2335_ _1607_ _1797_ VGND VGND VPWR VPWR _2632_ sky130_fd_sc_hd__nand4_1
XFILLER_0_10_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4184_ _0947_ _3143_ _3290_ VGND VGND VPWR VPWR _3291_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6825_ _2369_ _2370_ _2393_ _2394_ VGND VGND VPWR VPWR _2395_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3968_ net11 VGND VGND VPWR VPWR _2598_ sky130_fd_sc_hd__clkbuf_4
X_6756_ _0783_ _3156_ VGND VGND VPWR VPWR _2319_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5707_ _1168_ _1171_ VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__xnor2_2
X_3899_ _1788_ _1832_ _0936_ VGND VGND VPWR VPWR _1843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6687_ _1971_ _1973_ VGND VGND VPWR VPWR _2244_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5638_ _3343_ _0491_ _1094_ _1095_ VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__and4_1
XFILLER_0_60_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5569_ _1876_ _1008_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7308_ _2920_ _2921_ VGND VGND VPWR VPWR _2922_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7239_ _2845_ _2846_ _2804_ _2805_ VGND VGND VPWR VPWR _2848_ sky130_fd_sc_hd__o211a_1
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4940_ _0239_ _0244_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4871_ _0136_ _0137_ _0138_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_86_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6610_ _2157_ _2158_ VGND VGND VPWR VPWR _2159_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3822_ _0991_ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__buf_4
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6541_ _2070_ _2082_ _2083_ VGND VGND VPWR VPWR _2085_ sky130_fd_sc_hd__nand3_2
X_3753_ _0183_ _0226_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6472_ _1860_ _1866_ _1859_ VGND VGND VPWR VPWR _2009_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5423_ _2609_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__clkbuf_4
X_5354_ _3449_ _3448_ _2521_ _2565_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__nand4_2
XFILLER_0_11_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4305_ _0860_ _3410_ VGND VGND VPWR VPWR _3411_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5285_ _3056_ _0196_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__or2_1
X_4236_ _0324_ net60 _3313_ _3312_ VGND VGND VPWR VPWR _3342_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7024_ _2448_ _2449_ _2471_ _2472_ VGND VGND VPWR VPWR _2613_ sky130_fd_sc_hd__or4_1
X_4167_ _2456_ _3273_ VGND VGND VPWR VPWR _3274_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4098_ _3194_ _3199_ _3200_ _3201_ _3205_ VGND VGND VPWR VPWR _3206_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6808_ _0174_ _2784_ _2510_ _3720_ VGND VGND VPWR VPWR _2376_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6739_ _2007_ _2299_ VGND VGND VPWR VPWR _2300_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5070_ _2313_ _3619_ _0474_ _0475_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__nand4_2
X_4021_ _2609_ _1865_ _0892_ VGND VGND VPWR VPWR _3130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5972_ _0438_ _1451_ _1277_ VGND VGND VPWR VPWR _1462_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4923_ _0007_ _0306_ _0311_ _0316_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4854_ _2423_ net162 net31 VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4785_ _0163_ _0165_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__xnor2_1
X_3805_ _0150_ _0772_ _0805_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3736_ _0052_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6524_ _2401_ _1007_ VGND VGND VPWR VPWR _2066_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6455_ _1720_ _1851_ _1882_ _1883_ VGND VGND VPWR VPWR _1990_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_42_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5406_ _0849_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__buf_2
X_6386_ _1912_ _1913_ _1739_ _1814_ VGND VGND VPWR VPWR _1915_ sky130_fd_sc_hd__a211o_1
X_5337_ _0623_ _0642_ _0643_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__nand3_2
XFILLER_0_11_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5268_ _0692_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__clkbuf_2
X_4219_ _3240_ _3249_ _3248_ VGND VGND VPWR VPWR _3326_ sky130_fd_sc_hd__a21bo_1
X_7007_ _2375_ _2377_ _2592_ _2593_ VGND VGND VPWR VPWR _2594_ sky130_fd_sc_hd__o211ai_1
X_5199_ _3632_ _3633_ _3537_ _3651_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__and4_1
XFILLER_0_98_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4570_ _3670_ _3671_ _3517_ VGND VGND VPWR VPWR _3673_ sky130_fd_sc_hd__o21a_1
XFILLER_0_114_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6240_ _1625_ _1754_ _3305_ VGND VGND VPWR VPWR _1755_ sky130_fd_sc_hd__o21a_1
X_6171_ _1676_ _1677_ _1643_ _1644_ VGND VGND VPWR VPWR _1680_ sky130_fd_sc_hd__a211oi_2
X_5122_ _0530_ _0531_ _0400_ _0448_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__a211oi_2
X_5053_ _0451_ _0456_ _0457_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__and3_2
X_4004_ _0139_ _0772_ _0128_ VGND VGND VPWR VPWR _2991_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_79_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5955_ _1440_ _1442_ _1437_ VGND VGND VPWR VPWR _1444_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4906_ _0177_ _0180_ _0297_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5886_ _2117_ _0220_ VGND VGND VPWR VPWR _1368_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4837_ _0218_ _0221_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__xor2_2
XFILLER_0_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4768_ _0047_ _0056_ _0055_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_90_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4699_ _0069_ _0070_ _0016_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_120_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7487_ net96 net97 net98 _3113_ VGND VGND VPWR VPWR _3114_ sky130_fd_sc_hd__or4_1
X_6507_ _2030_ _2031_ _2046_ VGND VGND VPWR VPWR _2047_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6438_ _0346_ _0434_ net49 net50 VGND VGND VPWR VPWR _1971_ sky130_fd_sc_hd__and4_1
XFILLER_0_12_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6369_ _1894_ _1895_ VGND VGND VPWR VPWR _1896_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_8 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5740_ _3423_ _2248_ _3573_ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5671_ _1130_ _1131_ net130 net215 VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__a211oi_2
X_7410_ _3030_ _3033_ VGND VGND VPWR VPWR _3034_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4622_ _3709_ _3695_ _3723_ VGND VGND VPWR VPWR _3724_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4553_ _3536_ _3538_ _3539_ VGND VGND VPWR VPWR _3656_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_102_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7341_ _2793_ _2794_ VGND VGND VPWR VPWR _2959_ sky130_fd_sc_hd__or2b_1
XFILLER_0_52_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4484_ _3580_ _3583_ _3586_ _3587_ VGND VGND VPWR VPWR _3588_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7272_ _2880_ _2882_ VGND VGND VPWR VPWR _2883_ sky130_fd_sc_hd__nand2_2
XFILLER_0_111_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6223_ _1698_ _1699_ _1735_ _1736_ VGND VGND VPWR VPWR _1737_ sky130_fd_sc_hd__nor4_1
XFILLER_0_0_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6154_ _2160_ _0219_ _1524_ _1523_ _3719_ VGND VGND VPWR VPWR _1661_ sky130_fd_sc_hd__a32o_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5105_ _0511_ _0512_ _0513_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__a21o_1
X_6085_ net154 _1424_ _1584_ _1585_ VGND VGND VPWR VPWR _1586_ sky130_fd_sc_hd__a211o_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _0438_ _0439_ _0000_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6987_ _2456_ _2127_ _1169_ _1295_ VGND VGND VPWR VPWR _2572_ sky130_fd_sc_hd__and4_1
XFILLER_0_137_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5938_ _1357_ _1358_ _1422_ _1423_ VGND VGND VPWR VPWR _1425_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_63_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5869_ _1341_ _1348_ VGND VGND VPWR VPWR _1349_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_35_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput78 net78 VGND VGND VPWR VPWR result[18] sky130_fd_sc_hd__clkbuf_4
Xoutput89 net89 VGND VGND VPWR VPWR result[28] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_730 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6910_ _2485_ _2486_ _2327_ _2328_ VGND VGND VPWR VPWR _2488_ sky130_fd_sc_hd__a211o_1
XFILLER_0_134_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6841_ _2409_ _2410_ _2411_ VGND VGND VPWR VPWR _2413_ sky130_fd_sc_hd__or3b_2
XFILLER_0_134_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6772_ _0401_ net20 net21 _0499_ VGND VGND VPWR VPWR _2337_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3984_ net7 VGND VGND VPWR VPWR _2773_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5723_ _1186_ _1188_ net187 net118 VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_17_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5654_ _1110_ _1112_ _1113_ VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4605_ _3486_ _3707_ _3201_ VGND VGND VPWR VPWR _3708_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7324_ _3685_ _1876_ VGND VGND VPWR VPWR _2940_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_590 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5585_ _0335_ _0720_ _0873_ _0434_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4536_ _3630_ _3637_ _3638_ VGND VGND VPWR VPWR _3639_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4467_ _0652_ VGND VGND VPWR VPWR _3571_ sky130_fd_sc_hd__buf_4
X_7255_ _2863_ _2865_ _0320_ VGND VGND VPWR VPWR _2866_ sky130_fd_sc_hd__o21ai_1
X_6206_ _1563_ _1568_ _1562_ VGND VGND VPWR VPWR _1718_ sky130_fd_sc_hd__a21bo_1
X_4398_ _3108_ _3056_ _3200_ _3502_ VGND VGND VPWR VPWR _3503_ sky130_fd_sc_hd__a211o_1
X_7186_ _2718_ _0689_ VGND VGND VPWR VPWR _2790_ sky130_fd_sc_hd__nand2_1
X_6137_ _1418_ net109 _1579_ _1580_ VGND VGND VPWR VPWR _1642_ sky130_fd_sc_hd__o211a_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ _2881_ _2565_ VGND VGND VPWR VPWR _1567_ sky130_fd_sc_hd__nand2_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5019_ _3135_ _0328_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__nor2_1
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_395 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5370_ _0766_ _0767_ _0801_ _0802_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4321_ _1002_ _3425_ VGND VGND VPWR VPWR _3426_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4252_ _3242_ _3176_ net30 net31 VGND VGND VPWR VPWR _3358_ sky130_fd_sc_hd__nand4_2
XFILLER_0_10_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7040_ _2335_ _1607_ _1797_ _0117_ VGND VGND VPWR VPWR _2630_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4183_ _0947_ _3147_ VGND VGND VPWR VPWR _3290_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_468 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6824_ _2391_ _2392_ _2371_ _2372_ VGND VGND VPWR VPWR _2394_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_46_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3967_ _2576_ VGND VGND VPWR VPWR _2587_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6755_ _0854_ _2300_ _2317_ VGND VGND VPWR VPWR _2318_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5706_ _1002_ _1170_ VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3898_ _1810_ _1821_ _0892_ VGND VGND VPWR VPWR _1832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6686_ _2061_ _2069_ _2242_ VGND VGND VPWR VPWR _2243_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_143_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5637_ _3430_ _0491_ _1094_ _1095_ VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_5_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5568_ _0199_ _0848_ _1018_ _1019_ _0849_ VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__o311a_1
XFILLER_0_130_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4519_ _0477_ _3620_ _3617_ _3621_ VGND VGND VPWR VPWR _3622_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7307_ _2841_ _2843_ _1034_ _2299_ VGND VGND VPWR VPWR _2921_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5499_ _0942_ _0943_ _0923_ _0924_ VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__a211oi_2
X_7238_ _2804_ _2805_ _2845_ _2846_ VGND VGND VPWR VPWR _2847_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_111_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7169_ _2769_ _2770_ VGND VGND VPWR VPWR _2771_ sky130_fd_sc_hd__nor2_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4870_ _0255_ _0256_ _0254_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3821_ _0466_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6540_ _1836_ _1838_ _2081_ VGND VGND VPWR VPWR _2083_ sky130_fd_sc_hd__nand3_1
XFILLER_0_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3752_ _0183_ _0226_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6471_ _1999_ _2000_ _2005_ VGND VGND VPWR VPWR _2008_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5422_ _0848_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5353_ _0390_ _2521_ net10 _0488_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4304_ _3108_ _3210_ _3409_ _3200_ VGND VGND VPWR VPWR _3410_ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5284_ _3066_ _3500_ _0187_ _0710_ _0429_ _0189_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4235_ _3308_ VGND VGND VPWR VPWR _3341_ sky130_fd_sc_hd__inv_2
X_7023_ _2471_ VGND VGND VPWR VPWR _2612_ sky130_fd_sc_hd__inv_2
X_4166_ _3272_ VGND VGND VPWR VPWR _3273_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4097_ _1187_ _3202_ _3203_ _3204_ VGND VGND VPWR VPWR _3205_ sky130_fd_sc_hd__o22a_1
XFILLER_0_148_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6807_ _3720_ _0174_ _2784_ _2510_ VGND VGND VPWR VPWR _2375_ sky130_fd_sc_hd__and4_1
XFILLER_0_19_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4999_ _0356_ _0358_ _0396_ _0397_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__o22a_1
XFILLER_0_92_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6738_ net53 VGND VGND VPWR VPWR _2299_ sky130_fd_sc_hd__buf_2
XFILLER_0_34_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6669_ _2218_ _2223_ VGND VGND VPWR VPWR _2224_ sky130_fd_sc_hd__xor2_2
XFILLER_0_34_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_724 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4020_ _3128_ _2587_ _0903_ VGND VGND VPWR VPWR _3129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5971_ _3126_ _3285_ _3161_ VGND VGND VPWR VPWR _1461_ sky130_fd_sc_hd__a21o_1
XFILLER_0_149_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4922_ _3580_ _0312_ _0315_ _3587_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4853_ _2379_ _3430_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4784_ _3674_ _0164_ _0073_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3804_ _0150_ _0772_ _0794_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3735_ _0041_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__buf_6
XFILLER_0_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6523_ _2063_ _2064_ VGND VGND VPWR VPWR _2065_ sky130_fd_sc_hd__or2b_1
XFILLER_0_144_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_532 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6454_ _1848_ _1850_ _1910_ _1911_ VGND VGND VPWR VPWR _1989_ sky130_fd_sc_hd__nor4_1
X_5405_ _0575_ _0842_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6385_ _1739_ net105 _1912_ _1913_ VGND VGND VPWR VPWR _1914_ sky130_fd_sc_hd__o211ai_4
X_5336_ _0764_ _0765_ _0745_ _0746_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_11_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5267_ _0690_ _0691_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__or2_1
X_4218_ _3322_ _3323_ _3315_ VGND VGND VPWR VPWR _3325_ sky130_fd_sc_hd__a21o_1
X_7006_ _2664_ _0689_ _2590_ _2591_ VGND VGND VPWR VPWR _2593_ sky130_fd_sc_hd__nand4_2
XFILLER_0_98_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5198_ _3271_ _2204_ _2248_ _3632_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__a22oi_1
X_4149_ _3186_ _3231_ net159 _3256_ VGND VGND VPWR VPWR _3257_ sky130_fd_sc_hd__a211o_1
XFILLER_0_97_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire104 net200 VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_53_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6170_ _1643_ _1644_ _1676_ _1677_ VGND VGND VPWR VPWR _1678_ sky130_fd_sc_hd__o211a_1
X_5121_ _0400_ _0448_ _0530_ _0531_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__o211a_2
XFILLER_0_110_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5052_ _0445_ _0991_ _0327_ _0454_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__nand4_1
XFILLER_0_46_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4003_ _0794_ VGND VGND VPWR VPWR _2980_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5954_ net206 _1440_ _1442_ VGND VGND VPWR VPWR _1443_ sky130_fd_sc_hd__nand3_1
XFILLER_0_87_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4905_ _0174_ _3133_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__and2b_1
X_5885_ _1365_ _1366_ VGND VGND VPWR VPWR _1367_ sky130_fd_sc_hd__or2b_1
XFILLER_0_48_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4836_ _0466_ _0220_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4767_ _0143_ _0144_ _0135_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6506_ _2036_ _2045_ VGND VGND VPWR VPWR _2046_ sky130_fd_sc_hd__xor2_2
XFILLER_0_43_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4698_ _0016_ _0069_ _0070_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__or3_4
XFILLER_0_113_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7486_ net95 net80 net94 net91 VGND VGND VPWR VPWR _3113_ sky130_fd_sc_hd__or4_4
XFILLER_0_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6437_ _0357_ net48 _1817_ _1816_ VGND VGND VPWR VPWR _1970_ sky130_fd_sc_hd__a31o_1
XFILLER_0_101_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6368_ _0105_ _2773_ _2489_ _0104_ VGND VGND VPWR VPWR _1895_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5319_ _0614_ _0622_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__or2b_1
XFILLER_0_87_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6299_ _0357_ net48 VGND VGND VPWR VPWR _1819_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_9 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5670_ net130 net215 _1130_ _1131_ VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__o211a_4
XFILLER_0_85_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4621_ _3721_ _3722_ VGND VGND VPWR VPWR _3723_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4552_ _3652_ _3653_ _3650_ VGND VGND VPWR VPWR _3655_ sky130_fd_sc_hd__a21o_1
X_7340_ _2237_ _1170_ VGND VGND VPWR VPWR _2957_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4483_ _1701_ VGND VGND VPWR VPWR _3587_ sky130_fd_sc_hd__clkbuf_4
X_7271_ _0571_ net57 VGND VGND VPWR VPWR _2882_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6222_ _1732_ _1733_ _1573_ _1700_ VGND VGND VPWR VPWR _1736_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6153_ _1502_ _1505_ VGND VGND VPWR VPWR _1660_ sky130_fd_sc_hd__nand2_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5104_ _0511_ _0512_ _0513_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__nand3_2
X_6084_ _1518_ _1519_ _1582_ _1583_ VGND VGND VPWR VPWR _1585_ sky130_fd_sc_hd__a22oi_2
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _3135_ _0328_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__nand2_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6986_ _2570_ VGND VGND VPWR VPWR _2571_ sky130_fd_sc_hd__inv_2
X_5937_ _1357_ _1358_ _1422_ _1423_ VGND VGND VPWR VPWR _1424_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_48_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5868_ _1346_ _1347_ VGND VGND VPWR VPWR _1348_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4819_ _3580_ _0200_ _0202_ _3587_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__o211a_1
X_5799_ _1008_ _1876_ VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__and2b_1
XFILLER_0_105_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7469_ _1701_ _3085_ _3095_ VGND VGND VPWR VPWR _3096_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_31_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput79 net79 VGND VGND VPWR VPWR result[19] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6840_ _2205_ _2207_ _2203_ VGND VGND VPWR VPWR _2411_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_147_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6771_ _0881_ _0521_ net20 net21 VGND VGND VPWR VPWR _2336_ sky130_fd_sc_hd__nand4_2
XFILLER_0_57_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3983_ _2751_ VGND VGND VPWR VPWR _2762_ sky130_fd_sc_hd__buf_4
X_5722_ net187 net118 _1186_ _1188_ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5653_ _1110_ _1112_ _1113_ VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__nand3_1
XFILLER_0_73_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5584_ _0923_ _0924_ _0942_ _0943_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_72_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4604_ _3046_ _3591_ _3490_ VGND VGND VPWR VPWR _3707_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4535_ _1275_ _3631_ _3634_ _3636_ VGND VGND VPWR VPWR _3638_ sky130_fd_sc_hd__a22o_1
X_7323_ _3198_ _1778_ VGND VGND VPWR VPWR _2939_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4466_ _3479_ _3568_ _3305_ VGND VGND VPWR VPWR _3570_ sky130_fd_sc_hd__o21a_1
X_7254_ _2864_ _2662_ _2497_ _2663_ VGND VGND VPWR VPWR _2865_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_41_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6205_ _1708_ _1709_ _1715_ VGND VGND VPWR VPWR _1717_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4397_ _3108_ _3501_ VGND VGND VPWR VPWR _3502_ sky130_fd_sc_hd__nor2_1
X_7185_ _0420_ _2788_ VGND VGND VPWR VPWR _2789_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6136_ _1639_ _1640_ VGND VGND VPWR VPWR _1641_ sky130_fd_sc_hd__nor2_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6067_ _1854_ _1564_ _1565_ VGND VGND VPWR VPWR _1566_ sky130_fd_sc_hd__a21bo_1
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5018_ _2784_ _0327_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__and2_2
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6969_ _3620_ _2543_ _2383_ _2382_ _2609_ VGND VGND VPWR VPWR _2552_ sky130_fd_sc_hd__a32o_1
XFILLER_0_36_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4320_ _3424_ VGND VGND VPWR VPWR _3425_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4251_ net55 net29 VGND VGND VPWR VPWR _3357_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4182_ _0838_ _3126_ _3285_ _3287_ _3288_ VGND VGND VPWR VPWR _3289_ sky130_fd_sc_hd__a311o_1
XFILLER_0_38_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6823_ _2371_ _2372_ _2391_ _2392_ VGND VGND VPWR VPWR _2393_ sky130_fd_sc_hd__a211o_2
XFILLER_0_148_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3966_ _2565_ VGND VGND VPWR VPWR _2576_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6754_ _0855_ _2301_ _2316_ _1277_ VGND VGND VPWR VPWR _2317_ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6685_ _2067_ _2068_ VGND VGND VPWR VPWR _2242_ sky130_fd_sc_hd__or2b_1
X_5705_ _1169_ VGND VGND VPWR VPWR _1170_ sky130_fd_sc_hd__buf_4
XFILLER_0_143_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3897_ net20 VGND VGND VPWR VPWR _1821_ sky130_fd_sc_hd__clkbuf_4
X_5636_ _3195_ _3431_ net5 net6 VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__nand4_1
XFILLER_0_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5567_ _0428_ _1122_ _0005_ _0189_ VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_5_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5498_ _0923_ _0924_ _0942_ _0943_ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__o211a_1
X_4518_ _3616_ VGND VGND VPWR VPWR _3621_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7306_ _1034_ _2299_ _2841_ _2843_ VGND VGND VPWR VPWR _2920_ sky130_fd_sc_hd__a211oi_1
X_4449_ _3550_ _3551_ _3462_ _3464_ VGND VGND VPWR VPWR _3553_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7237_ _2843_ _2844_ _2603_ _2605_ VGND VGND VPWR VPWR _2846_ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7168_ _2127_ _2171_ _1170_ _1295_ VGND VGND VPWR VPWR _2770_ sky130_fd_sc_hd__and4_1
X_6119_ _1437_ _1440_ _1597_ VGND VGND VPWR VPWR _1622_ sky130_fd_sc_hd__or3_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7099_ _2051_ net56 VGND VGND VPWR VPWR _2694_ sky130_fd_sc_hd__nor2_1
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3820_ _0303_ VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3751_ _0215_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__buf_4
XFILLER_0_125_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_703 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6470_ _1999_ _2000_ _2005_ VGND VGND VPWR VPWR _2006_ sky130_fd_sc_hd__nand3_1
XFILLER_0_40_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5421_ _0823_ _0825_ _0859_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__o21ai_4
XFILLER_0_70_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5352_ _0292_ net8 VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4303_ _3077_ _1089_ _3408_ _1723_ VGND VGND VPWR VPWR _3409_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5283_ _3128_ _0558_ _3135_ _3134_ _3046_ _0584_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__mux4_1
X_7022_ _2607_ _2608_ net213 _2440_ VGND VGND VPWR VPWR _2611_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4234_ _3306_ _3307_ _3308_ VGND VGND VPWR VPWR _3340_ sky130_fd_sc_hd__or3_2
X_4165_ _3271_ VGND VGND VPWR VPWR _3272_ sky130_fd_sc_hd__buf_6
XFILLER_0_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4096_ _1220_ VGND VGND VPWR VPWR _3204_ sky130_fd_sc_hd__buf_2
XFILLER_0_78_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6806_ _2153_ _2161_ VGND VGND VPWR VPWR _2374_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4998_ _0356_ _0358_ _0396_ _0397_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__nor4_2
XFILLER_0_92_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_664 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6737_ _2277_ _2284_ _2294_ _2298_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__nand4_4
XFILLER_0_45_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3949_ _2379_ VGND VGND VPWR VPWR _2390_ sky130_fd_sc_hd__buf_6
XFILLER_0_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6668_ _2221_ _2222_ VGND VGND VPWR VPWR _2223_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6599_ _2140_ _2141_ _2146_ VGND VGND VPWR VPWR _2147_ sky130_fd_sc_hd__nand3_1
X_5619_ _2390_ _0219_ _1073_ _1074_ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__nand4_2
XFILLER_0_104_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5970_ _1452_ _1457_ _0419_ VGND VGND VPWR VPWR _1459_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4921_ _3580_ _0313_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__nand2_1
X_4852_ _0131_ _0132_ _0133_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_87_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3803_ _0783_ _0641_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4783_ _0071_ _0072_ _3670_ _3672_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_62_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3734_ _0030_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__buf_8
XFILLER_0_16_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6522_ _2127_ _0721_ _0874_ _2445_ VGND VGND VPWR VPWR _2064_ sky130_fd_sc_hd__a22o_1
X_6453_ _1986_ _1987_ VGND VGND VPWR VPWR _1988_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5404_ _0571_ _0840_ _0841_ _0839_ _0573_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6384_ _1848_ _1850_ _1910_ _1911_ VGND VGND VPWR VPWR _1913_ sky130_fd_sc_hd__o22ai_4
X_5335_ _0745_ _0746_ _0764_ _0765_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5266_ _3128_ _0689_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4217_ _3315_ _3322_ _3323_ VGND VGND VPWR VPWR _3324_ sky130_fd_sc_hd__nand3_1
XFILLER_0_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7005_ _2664_ _0689_ _2590_ _2591_ VGND VGND VPWR VPWR _2592_ sky130_fd_sc_hd__a22o_1
X_5197_ _0502_ _0503_ _0504_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__o21ba_1
X_4148_ _3253_ _3254_ _3235_ VGND VGND VPWR VPWR _3256_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4079_ _3186_ _3187_ VGND VGND VPWR VPWR _3188_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_807 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5120_ _0528_ _0529_ _0464_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5051_ _0445_ _0327_ _0454_ _0477_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4002_ _2936_ _2958_ VGND VGND VPWR VPWR _2969_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5953_ _1146_ _1149_ _1441_ VGND VGND VPWR VPWR _1442_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5884_ _2204_ _3718_ _0099_ _0247_ VGND VGND VPWR VPWR _1366_ sky130_fd_sc_hd__a22o_1
X_4904_ _0294_ _0295_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4835_ _0219_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_16_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4766_ _0135_ _0143_ _0144_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__nand3_1
XFILLER_0_90_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6505_ _2043_ _2044_ VGND VGND VPWR VPWR _2045_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4697_ _0067_ _0068_ _0017_ _3668_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_70_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7485_ net86 net87 net89 VGND VGND VPWR VPWR _3112_ sky130_fd_sc_hd__or3_4
XFILLER_0_113_363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6436_ _1820_ _1828_ _1826_ VGND VGND VPWR VPWR _1969_ sky130_fd_sc_hd__o21ai_1
X_6367_ _3423_ _0105_ _2773_ _2499_ VGND VGND VPWR VPWR _1894_ sky130_fd_sc_hd__nand4_1
X_5318_ _0615_ _0618_ _0620_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__or3_1
XFILLER_0_87_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6298_ _1816_ _1817_ VGND VGND VPWR VPWR _1818_ sky130_fd_sc_hd__or2b_1
X_5249_ _0650_ _0651_ _0670_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_97_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_636 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_670 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_523 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4620_ _2653_ _3718_ VGND VGND VPWR VPWR _3722_ sky130_fd_sc_hd__and2_2
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4551_ _3650_ _3652_ _3653_ VGND VGND VPWR VPWR _3654_ sky130_fd_sc_hd__nand3_1
XFILLER_0_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4482_ _3580_ _3585_ VGND VGND VPWR VPWR _3586_ sky130_fd_sc_hd__nand2_1
X_7270_ _0571_ net57 VGND VGND VPWR VPWR _2880_ sky130_fd_sc_hd__or2_1
X_6221_ _1573_ _1700_ _1732_ _1733_ VGND VGND VPWR VPWR _1735_ sky130_fd_sc_hd__o211a_2
XFILLER_0_0_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _1650_ _1658_ VGND VGND VPWR VPWR _1659_ sky130_fd_sc_hd__xor2_2
XFILLER_0_148_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5103_ _0378_ _0381_ _0382_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_110_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _1518_ _1519_ _1582_ _1583_ VGND VGND VPWR VPWR _1584_ sky130_fd_sc_hd__and4_2
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ net124 VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__clkbuf_4
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6985_ _2127_ _1169_ _1294_ _2456_ VGND VGND VPWR VPWR _2570_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5936_ net203 _1421_ _1249_ _1359_ VGND VGND VPWR VPWR _1423_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_48_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5867_ _1344_ _1345_ _1197_ _1200_ VGND VGND VPWR VPWR _1347_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4818_ _3580_ _0201_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5798_ _1270_ _1271_ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__nand2_4
XFILLER_0_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4749_ _3530_ _0035_ _0125_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_50_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7468_ _1646_ _3086_ _3090_ _3094_ VGND VGND VPWR VPWR _3095_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6419_ _1810_ _1949_ VGND VGND VPWR VPWR _1950_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7399_ _2931_ _3021_ VGND VGND VPWR VPWR _3022_ sky130_fd_sc_hd__xnor2_1
Xoutput69 net69 VGND VGND VPWR VPWR result[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3982_ _2740_ VGND VGND VPWR VPWR _2751_ sky130_fd_sc_hd__buf_6
X_6770_ _2151_ _2152_ _2162_ VGND VGND VPWR VPWR _2334_ sky130_fd_sc_hd__nor3_1
XFILLER_0_9_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5721_ _1184_ _1185_ _1172_ VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5652_ _0963_ _0964_ _0965_ VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_84_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4603_ _0860_ _3705_ VGND VGND VPWR VPWR _3706_ sky130_fd_sc_hd__nor2_1
X_5583_ _0905_ _0917_ _1036_ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4534_ _0205_ _3631_ _3634_ _3636_ VGND VGND VPWR VPWR _3637_ sky130_fd_sc_hd__nand4_2
X_7322_ _2826_ _2831_ _2832_ _2834_ _2825_ VGND VGND VPWR VPWR _2938_ sky130_fd_sc_hd__a32o_1
XFILLER_0_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4465_ _3479_ _3568_ VGND VGND VPWR VPWR _3569_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7253_ _2487_ _2500_ VGND VGND VPWR VPWR _2864_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6204_ _1708_ _1709_ _1715_ VGND VGND VPWR VPWR _1716_ sky130_fd_sc_hd__nand3_1
X_4396_ _3066_ _3500_ _3077_ VGND VGND VPWR VPWR _3501_ sky130_fd_sc_hd__mux2_1
X_7184_ _2762_ _0454_ VGND VGND VPWR VPWR _2788_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6135_ _1516_ _1518_ _1638_ VGND VGND VPWR VPWR _1640_ sky130_fd_sc_hd__and3_1
X_6066_ _0030_ net11 net13 _3169_ VGND VGND VPWR VPWR _1565_ sky130_fd_sc_hd__a22o_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5017_ _2980_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__clkbuf_4
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6968_ _3685_ _2576_ _2548_ _2549_ VGND VGND VPWR VPWR _2551_ sky130_fd_sc_hd__nand4_4
XFILLER_0_49_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5919_ _1401_ _1402_ _1403_ VGND VGND VPWR VPWR _1404_ sky130_fd_sc_hd__nand3_1
XFILLER_0_91_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6899_ _2475_ VGND VGND VPWR VPWR _2476_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_816 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4250_ _3351_ _3355_ VGND VGND VPWR VPWR _3356_ sky130_fd_sc_hd__xor2_2
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4181_ net123 _3274_ _3275_ _1187_ _3162_ VGND VGND VPWR VPWR _3288_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6822_ _2373_ _2374_ _2389_ VGND VGND VPWR VPWR _2392_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_662 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3965_ net10 VGND VGND VPWR VPWR _2565_ sky130_fd_sc_hd__buf_4
XFILLER_0_70_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6753_ _3589_ _2300_ _2301_ VGND VGND VPWR VPWR _2316_ sky130_fd_sc_hd__o21ai_1
X_3896_ _1799_ VGND VGND VPWR VPWR _1810_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6684_ _2087_ _2089_ VGND VGND VPWR VPWR _2241_ sky130_fd_sc_hd__nand2_1
X_5704_ net46 VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__clkbuf_4
X_5635_ net162 net5 net6 _3433_ VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5566_ _0585_ _1017_ _0429_ VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5497_ _0926_ _0927_ _0941_ VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__nand3_2
X_4517_ _3619_ VGND VGND VPWR VPWR _3620_ sky130_fd_sc_hd__buf_4
X_7305_ _2917_ _2918_ VGND VGND VPWR VPWR _2919_ sky130_fd_sc_hd__nor2_1
X_4448_ _3462_ _3464_ _3550_ _3551_ VGND VGND VPWR VPWR _3552_ sky130_fd_sc_hd__a211o_4
X_7236_ _2603_ _2605_ _2843_ _2844_ VGND VGND VPWR VPWR _2845_ sky130_fd_sc_hd__a211oi_4
X_4379_ _3482_ _3483_ VGND VGND VPWR VPWR _3484_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7167_ _2171_ _1170_ _1295_ _2127_ VGND VGND VPWR VPWR _2769_ sky130_fd_sc_hd__a22oi_1
X_6118_ _1597_ _1598_ VGND VGND VPWR VPWR _1621_ sky130_fd_sc_hd__or2_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7098_ _2693_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_1
X_6049_ _3632_ _3633_ _2489_ _2521_ VGND VGND VPWR VPWR _1546_ sky130_fd_sc_hd__nand4_2
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3750_ _0205_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5420_ _0181_ _0832_ _0833_ _0837_ _0858_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__o311a_2
XFILLER_0_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5351_ _0779_ _0782_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__xor2_2
XFILLER_0_2_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4302_ _3077_ _3407_ VGND VGND VPWR VPWR _3408_ sky130_fd_sc_hd__nand2_1
X_5282_ _0704_ _0705_ _0706_ _3161_ _0708_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4233_ _3279_ _3280_ _3304_ _3339_ VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__a211o_4
X_7021_ net213 _2440_ _2607_ _2608_ VGND VGND VPWR VPWR _2610_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4164_ _3270_ VGND VGND VPWR VPWR _3271_ sky130_fd_sc_hd__clkbuf_4
X_4095_ _1209_ _3199_ _3202_ VGND VGND VPWR VPWR _3203_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6805_ _2154_ _2159_ VGND VGND VPWR VPWR _2373_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4997_ _0394_ _0395_ _0266_ _0359_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__o211a_1
X_6736_ _2280_ _2296_ _2297_ VGND VGND VPWR VPWR _2298_ sky130_fd_sc_hd__o21ai_1
X_3948_ _2368_ VGND VGND VPWR VPWR _2379_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3879_ _0183_ _1384_ _1395_ VGND VGND VPWR VPWR _1624_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6667_ _2226_ _0688_ _2219_ _2220_ VGND VGND VPWR VPWR _2222_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_60_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6598_ _2144_ _2145_ VGND VGND VPWR VPWR _2146_ sky130_fd_sc_hd__xor2_1
X_5618_ _2390_ _0220_ _1073_ _1074_ VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5549_ _0722_ _2587_ VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__and2b_1
XFILLER_0_42_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7219_ _2572_ _2574_ VGND VGND VPWR VPWR _2826_ sky130_fd_sc_hd__or2_1
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4920_ _0196_ _2062_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__or2b_1
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4851_ _2324_ _3385_ _0125_ _0035_ _2445_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__a32o_1
XFILLER_0_59_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3802_ net65 VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4782_ _0160_ _0162_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_16_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3733_ net59 VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__buf_8
XFILLER_0_82_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6521_ _2445_ _2127_ _0721_ _0874_ VGND VGND VPWR VPWR _2063_ sky130_fd_sc_hd__and4_1
XFILLER_0_141_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6452_ _1807_ _1634_ _1805_ VGND VGND VPWR VPWR _1987_ sky130_fd_sc_hd__and3b_1
XFILLER_0_43_646 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5403_ _0199_ _3727_ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_578 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6383_ _1848_ _1850_ _1910_ _1911_ VGND VGND VPWR VPWR _1912_ sky130_fd_sc_hd__or4_4
X_5334_ _0747_ _0748_ _0763_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__nand3_2
X_5265_ _3128_ _0689_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__and2_1
X_4216_ _3319_ _3320_ _3321_ VGND VGND VPWR VPWR _3323_ sky130_fd_sc_hd__a21o_1
X_5196_ _3388_ _0493_ _0494_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__a21boi_2
X_7004_ _2718_ _2762_ _0328_ _0559_ VGND VGND VPWR VPWR _2591_ sky130_fd_sc_hd__nand4_2
XFILLER_0_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4147_ _3235_ _3253_ _3254_ VGND VGND VPWR VPWR _3255_ sky130_fd_sc_hd__nor3_2
X_4078_ _3168_ _1515_ _3185_ VGND VGND VPWR VPWR _3187_ sky130_fd_sc_hd__or3_4
XFILLER_0_97_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire106 _0986_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__buf_2
XFILLER_0_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6719_ _1821_ _2263_ VGND VGND VPWR VPWR _2279_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5050_ _0453_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__clkbuf_4
X_4001_ _0150_ _0608_ _2947_ VGND VGND VPWR VPWR _2958_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5952_ _1142_ _1267_ VGND VGND VPWR VPWR _1441_ sky130_fd_sc_hd__or2_1
X_4903_ _2762_ _0293_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__nand2_2
XFILLER_0_62_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5883_ _0247_ _2204_ _3718_ _0099_ VGND VGND VPWR VPWR _1365_ sky130_fd_sc_hd__and4_1
XFILLER_0_62_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4834_ net38 VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4765_ _0140_ _0141_ _0142_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6504_ _2039_ _2041_ _2042_ VGND VGND VPWR VPWR _2044_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_71_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4696_ _0017_ _3668_ _0067_ _0068_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7484_ _3587_ _3099_ _3105_ _3111_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__a211o_1
XFILLER_0_71_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6435_ _1846_ _1848_ VGND VGND VPWR VPWR _1968_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6366_ _1891_ _1892_ VGND VGND VPWR VPWR _1893_ sky130_fd_sc_hd__nand2_1
X_5317_ _0599_ _0606_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6297_ _0106_ net46 net47 _0205_ VGND VGND VPWR VPWR _1817_ sky130_fd_sc_hd__a22o_1
X_5248_ _0650_ _0651_ _0670_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__nor3b_4
X_5179_ _3440_ _3635_ _0340_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4550_ _3451_ _3452_ _3537_ _3651_ VGND VGND VPWR VPWR _3653_ sky130_fd_sc_hd__nand4_2
XFILLER_0_106_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4481_ _3301_ _3584_ VGND VGND VPWR VPWR _3585_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6220_ _1720_ _1721_ _1731_ VGND VGND VPWR VPWR _1733_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6151_ _1655_ _1656_ VGND VGND VPWR VPWR _1658_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5102_ _0508_ _0509_ _0507_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6082_ _1579_ _1580_ _1418_ net109 VGND VGND VPWR VPWR _1583_ sky130_fd_sc_hd__a211o_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _3194_ _0420_ _0421_ _3414_ _3201_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__a221o_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6984_ _2373_ _2374_ _2389_ VGND VGND VPWR VPWR _2569_ sky130_fd_sc_hd__a21o_1
X_5935_ _1249_ _1359_ net203 _1421_ VGND VGND VPWR VPWR _1422_ sky130_fd_sc_hd__a211o_1
XFILLER_0_91_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5866_ _1197_ _1200_ _1344_ _1345_ VGND VGND VPWR VPWR _1346_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4817_ _3490_ _3486_ _3145_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5797_ _1909_ _1170_ VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__nand2_2
XFILLER_0_16_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4748_ _3195_ _2423_ _3633_ _2368_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4679_ _3449_ _3448_ _3651_ _2642_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__nand4_2
XFILLER_0_102_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7467_ _3091_ _3265_ _3092_ _3093_ _3595_ VGND VGND VPWR VPWR _3094_ sky130_fd_sc_hd__o32a_1
XFILLER_0_31_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6418_ net51 VGND VGND VPWR VPWR _1949_ sky130_fd_sc_hd__buf_2
X_7398_ _2937_ _3020_ VGND VGND VPWR VPWR _3021_ sky130_fd_sc_hd__xnor2_1
X_6349_ _3433_ net162 net10 net11 VGND VGND VPWR VPWR _1874_ sky130_fd_sc_hd__and4_1
XFILLER_0_11_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3981_ net6 VGND VGND VPWR VPWR _2740_ sky130_fd_sc_hd__buf_4
XFILLER_0_69_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5720_ _1172_ _1184_ _1185_ VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__nand3_2
XFILLER_0_9_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5651_ _1108_ _1109_ _1107_ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5582_ _0915_ _0916_ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__and2b_1
X_4602_ _3486_ _3703_ _3704_ VGND VGND VPWR VPWR _3705_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_142_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4533_ _3440_ _3635_ _3632_ _3271_ VGND VGND VPWR VPWR _3636_ sky130_fd_sc_hd__nand4_2
X_7321_ _2932_ _2935_ VGND VGND VPWR VPWR _2937_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7252_ _2860_ _2862_ VGND VGND VPWR VPWR _2863_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_755 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4464_ _3566_ _3567_ VGND VGND VPWR VPWR _3568_ sky130_fd_sc_hd__or2_1
X_6203_ _1713_ _1714_ VGND VGND VPWR VPWR _1715_ sky130_fd_sc_hd__xor2_1
XFILLER_0_68_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7183_ _2543_ _2542_ _2545_ _2546_ VGND VGND VPWR VPWR _2787_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_68_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4395_ _2182_ _2138_ _3139_ _2412_ _0914_ _3131_ VGND VGND VPWR VPWR _3500_ sky130_fd_sc_hd__mux4_2
XFILLER_0_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6134_ _1516_ _1518_ _1638_ VGND VGND VPWR VPWR _1639_ sky130_fd_sc_hd__a21oi_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _3169_ net191 net11 VGND VGND VPWR VPWR _1564_ sky130_fd_sc_hd__and3_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ net209 _0417_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__xnor2_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6967_ _3685_ _2576_ _2548_ _2549_ VGND VGND VPWR VPWR _2550_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5918_ _0281_ net13 VGND VGND VPWR VPWR _1403_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6898_ _2231_ _2233_ _2473_ _2474_ VGND VGND VPWR VPWR _2475_ sky130_fd_sc_hd__a211o_1
XFILLER_0_134_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5849_ _0707_ _0477_ _1169_ _1294_ VGND VGND VPWR VPWR _1327_ sky130_fd_sc_hd__and4_1
XFILLER_0_17_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4180_ _3275_ _3286_ VGND VGND VPWR VPWR _3287_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6821_ _2373_ _2374_ _2389_ VGND VGND VPWR VPWR _2391_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_148_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3964_ _2510_ _2543_ _2029_ VGND VGND VPWR VPWR _2554_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_674 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6752_ _0003_ _0005_ _1018_ _2314_ _0867_ _0573_ VGND VGND VPWR VPWR _2315_ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3895_ net19 VGND VGND VPWR VPWR _1799_ sky130_fd_sc_hd__buf_2
X_5703_ _1166_ _1167_ VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6683_ _2238_ _2239_ VGND VGND VPWR VPWR _2240_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5634_ _2892_ _2751_ _0960_ _0959_ _2499_ VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__a32o_1
XFILLER_0_73_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5565_ _1876_ _0862_ _2587_ _3128_ _0583_ _0584_ VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7304_ _1023_ _2263_ _2845_ _2847_ VGND VGND VPWR VPWR _2918_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_41_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5496_ _0926_ _0927_ _0941_ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__a21o_2
X_4516_ net35 VGND VGND VPWR VPWR _3619_ sky130_fd_sc_hd__buf_2
X_4447_ _3548_ _3549_ net131 VGND VGND VPWR VPWR _3551_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7235_ _2841_ _2842_ _2821_ VGND VGND VPWR VPWR _2844_ sky130_fd_sc_hd__o21a_1
X_7166_ _2558_ _2560_ VGND VGND VPWR VPWR _2768_ sky130_fd_sc_hd__and2b_1
X_6117_ _1149_ _1618_ VGND VGND VPWR VPWR _1620_ sky130_fd_sc_hd__or2_4
X_4378_ _3387_ _3397_ _3388_ VGND VGND VPWR VPWR _3483_ sky130_fd_sc_hd__o21ba_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7097_ _2669_ _2676_ _2692_ VGND VGND VPWR VPWR _2693_ sky130_fd_sc_hd__or3b_1
X_6048_ _2881_ _2532_ _1397_ _1396_ _2598_ VGND VGND VPWR VPWR _1545_ sky130_fd_sc_hd__a32o_1
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_474 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_703 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5350_ _2773_ _0780_ _0781_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_2_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4301_ _2138_ _3139_ _2412_ _2346_ _0914_ _3131_ VGND VGND VPWR VPWR _3407_ sky130_fd_sc_hd__mux4_2
X_5281_ _3194_ _0690_ _0691_ _3414_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__a22o_1
X_4232_ _3305_ _3337_ _3338_ VGND VGND VPWR VPWR _3339_ sky130_fd_sc_hd__and3_1
X_7020_ _2564_ _2566_ _2605_ _2606_ VGND VGND VPWR VPWR _2608_ sky130_fd_sc_hd__a2bb2o_1
X_4163_ net62 VGND VGND VPWR VPWR _3270_ sky130_fd_sc_hd__buf_6
X_4094_ _2401_ _3198_ VGND VGND VPWR VPWR _3202_ sky130_fd_sc_hd__or2_2
XFILLER_0_148_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4996_ _0266_ _0359_ _0394_ _0395_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__a211oi_2
X_6804_ _2175_ _2183_ VGND VGND VPWR VPWR _2372_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3947_ net29 VGND VGND VPWR VPWR _2368_ sky130_fd_sc_hd__buf_4
XFILLER_0_46_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6735_ _2280_ _2296_ _0181_ VGND VGND VPWR VPWR _2297_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3878_ _1592_ _1603_ VGND VGND VPWR VPWR _1613_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6666_ _2219_ _2220_ _2226_ _0688_ VGND VGND VPWR VPWR _2221_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_143_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6597_ _2892_ _1931_ VGND VGND VPWR VPWR _2145_ sky130_fd_sc_hd__nand2_1
X_5617_ _2434_ _3644_ _0339_ _0340_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__nand4_4
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5548_ _0824_ _0997_ _0895_ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__or3_1
XFILLER_0_60_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5479_ _0760_ _0759_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__and2b_1
X_7218_ _1023_ _2346_ _1608_ _1797_ _2634_ VGND VGND VPWR VPWR _2825_ sky130_fd_sc_hd__a41o_1
X_7149_ _3513_ _1865_ _1898_ _3425_ VGND VGND VPWR VPWR _2749_ sky130_fd_sc_hd__a22oi_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4850_ _0130_ _0148_ _0149_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__nand3_1
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3801_ _0674_ _0761_ _0237_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__o21a_1
XFILLER_0_68_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4781_ _0069_ _0071_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__or2b_1
XFILLER_0_117_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6520_ _2059_ _2060_ VGND VGND VPWR VPWR _2061_ sky130_fd_sc_hd__nand2_2
XFILLER_0_15_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6451_ _1968_ _1984_ VGND VGND VPWR VPWR _1986_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6382_ _1907_ _1908_ _1735_ net201 VGND VGND VPWR VPWR _1911_ sky130_fd_sc_hd__a211oi_4
X_5402_ _3727_ _3707_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5333_ _0747_ _0748_ _0763_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__a21o_2
XFILLER_0_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5264_ _0688_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__clkbuf_4
X_5195_ _0501_ _0519_ _0520_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__nand3_2
X_4215_ _3319_ _3320_ _3321_ VGND VGND VPWR VPWR _3322_ sky130_fd_sc_hd__nand3_1
XFILLER_0_76_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7003_ _2762_ _0328_ _0559_ _2718_ VGND VGND VPWR VPWR _2590_ sky130_fd_sc_hd__a22o_1
X_4146_ _3250_ _3251_ _3252_ VGND VGND VPWR VPWR _3254_ sky130_fd_sc_hd__a21oi_1
X_4077_ _3168_ _1515_ _3185_ VGND VGND VPWR VPWR _3186_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4979_ _0372_ _0376_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__xor2_2
XFILLER_0_93_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6718_ _1821_ _2263_ VGND VGND VPWR VPWR _2278_ sky130_fd_sc_hd__or2_2
XFILLER_0_132_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6649_ _2200_ _2201_ VGND VGND VPWR VPWR _2202_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_786 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4000_ _0838_ _0117_ VGND VGND VPWR VPWR _2947_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5951_ _1265_ _1438_ _1267_ _1155_ VGND VGND VPWR VPWR _1440_ sky130_fd_sc_hd__o22a_1
XFILLER_0_153_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4902_ _3134_ _0293_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5882_ _1217_ _1225_ VGND VGND VPWR VPWR _1364_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4833_ _0216_ _0217_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4764_ _0140_ _0141_ _0142_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__nand3_1
XFILLER_0_117_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7483_ _1613_ _3106_ _3110_ VGND VGND VPWR VPWR _3111_ sky130_fd_sc_hd__o21ai_1
X_6503_ _2039_ _2041_ _2042_ VGND VGND VPWR VPWR _2043_ sky130_fd_sc_hd__or3b_4
XFILLER_0_71_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4695_ _0065_ _0066_ _0029_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6434_ _1475_ _1637_ _1812_ VGND VGND VPWR VPWR _1967_ sky130_fd_sc_hd__and3_1
XFILLER_0_141_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6365_ _2259_ _0220_ _1889_ _1890_ VGND VGND VPWR VPWR _1892_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5316_ _0605_ _0604_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6296_ _0095_ _0205_ net46 net47 VGND VGND VPWR VPWR _1816_ sky130_fd_sc_hd__and4_1
X_5247_ _0461_ _0669_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__xor2_1
X_5178_ _0215_ _0219_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4129_ net58 net59 _1264_ _0314_ VGND VGND VPWR VPWR _3237_ sky130_fd_sc_hd__and4_1
XFILLER_0_97_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4480_ _2062_ _3024_ _3224_ _3077_ VGND VGND VPWR VPWR _3584_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6150_ _1489_ _1491_ VGND VGND VPWR VPWR _1656_ sky130_fd_sc_hd__or2_1
X_5101_ _0507_ _0508_ _0509_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__nand3_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _1418_ net109 _1579_ _1580_ VGND VGND VPWR VPWR _1582_ sky130_fd_sc_hd__o211ai_2
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _3285_ _0435_ _0189_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__mux2_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6983_ _2418_ _2431_ _2432_ VGND VGND VPWR VPWR _2568_ sky130_fd_sc_hd__and3_1
X_5934_ _1381_ _1382_ _1418_ _1419_ VGND VGND VPWR VPWR _1421_ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5865_ _2313_ _0654_ _1342_ _1343_ VGND VGND VPWR VPWR _1345_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_48_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4816_ _3132_ _3136_ _3148_ _3151_ _3087_ _0199_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__mux4_1
XFILLER_0_29_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5796_ _1909_ _1170_ VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__or2_2
XFILLER_0_133_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4747_ _2313_ _3631_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4678_ _0390_ _3651_ _2642_ _0488_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__a22o_1
X_7466_ _0259_ _0761_ VGND VGND VPWR VPWR _3093_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6417_ _0320_ _1927_ _1934_ _1948_ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__a211o_2
X_7397_ _2938_ _3019_ VGND VGND VPWR VPWR _3020_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6348_ _2892_ _2598_ _1711_ _1710_ _1898_ VGND VGND VPWR VPWR _1873_ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6279_ net50 VGND VGND VPWR VPWR _1797_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3980_ _2675_ _2718_ _2029_ VGND VGND VPWR VPWR _2729_ sky130_fd_sc_hd__mux2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5650_ _1107_ _1108_ _1109_ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__nand3_1
XFILLER_0_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4601_ _3087_ _3284_ _3301_ VGND VGND VPWR VPWR _3704_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5581_ _0898_ _0899_ _0919_ _0920_ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__a211o_1
XFILLER_0_72_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4532_ net28 VGND VGND VPWR VPWR _3635_ sky130_fd_sc_hd__clkbuf_4
X_7320_ _2933_ _2934_ VGND VGND VPWR VPWR _2935_ sky130_fd_sc_hd__xor2_1
XFILLER_0_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4463_ _3564_ _3565_ _3476_ VGND VGND VPWR VPWR _3567_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7251_ _2660_ _2859_ VGND VGND VPWR VPWR _2862_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6202_ _2881_ _2598_ VGND VGND VPWR VPWR _1714_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4394_ _3482_ _3497_ _3498_ VGND VGND VPWR VPWR _3499_ sky130_fd_sc_hd__o21a_1
X_7182_ _2591_ _2593_ VGND VGND VPWR VPWR _2786_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6133_ _1475_ _1637_ VGND VGND VPWR VPWR _1638_ sky130_fd_sc_hd__xnor2_1
X_6064_ _1558_ _1560_ _1561_ VGND VGND VPWR VPWR _1563_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _0287_ _0289_ _0416_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__a21o_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6966_ _3424_ _3513_ _2609_ _1865_ VGND VGND VPWR VPWR _2549_ sky130_fd_sc_hd__nand4_4
X_5917_ net178 _1887_ net15 _3242_ VGND VGND VPWR VPWR _1402_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6897_ _2448_ _2449_ _2471_ _2472_ VGND VGND VPWR VPWR _2474_ sky130_fd_sc_hd__o22a_1
XFILLER_0_119_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5848_ _1325_ VGND VGND VPWR VPWR _1326_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_580 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5779_ _1215_ _1216_ _1249_ _1250_ VGND VGND VPWR VPWR _1251_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_17_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7449_ _0510_ _3210_ VGND VGND VPWR VPWR _3075_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6820_ _2381_ _2388_ VGND VGND VPWR VPWR _2389_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3963_ _2532_ VGND VGND VPWR VPWR _2543_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6751_ _1758_ _2312_ _0866_ VGND VGND VPWR VPWR _2314_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3894_ _1756_ _1778_ _0892_ VGND VGND VPWR VPWR _1788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6682_ _2054_ _2091_ VGND VGND VPWR VPWR _2239_ sky130_fd_sc_hd__and2b_1
X_5702_ _1041_ _1042_ _1040_ VGND VGND VPWR VPWR _1167_ sky130_fd_sc_hd__o21ai_2
X_5633_ _3197_ _3272_ _2664_ _2707_ _0953_ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__a41o_1
XFILLER_0_26_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5564_ _1011_ _1014_ _0181_ VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4515_ _3616_ net35 net1 _3617_ VGND VGND VPWR VPWR _3618_ sky130_fd_sc_hd__and4b_1
XFILLER_0_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7303_ _2845_ _2847_ _1023_ _2263_ VGND VGND VPWR VPWR _2917_ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5495_ _0932_ _0940_ VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__xnor2_2
X_4446_ net131 _3548_ _3549_ VGND VGND VPWR VPWR _3550_ sky130_fd_sc_hd__and3_1
X_7234_ _2821_ _2841_ _2842_ VGND VGND VPWR VPWR _2843_ sky130_fd_sc_hd__nor3_2
X_4377_ _3480_ _3481_ VGND VGND VPWR VPWR _3482_ sky130_fd_sc_hd__or2_2
X_7165_ _2586_ _2600_ _2599_ VGND VGND VPWR VPWR _2767_ sky130_fd_sc_hd__a21bo_1
X_6116_ _0549_ _0552_ _0553_ _1145_ _1618_ VGND VGND VPWR VPWR _1619_ sky130_fd_sc_hd__a311o_4
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7096_ _2678_ _2679_ _2691_ VGND VGND VPWR VPWR _2692_ sky130_fd_sc_hd__a21oi_1
X_6047_ _1387_ _1389_ VGND VGND VPWR VPWR _1544_ sky130_fd_sc_hd__nand2_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6949_ _2528_ _2529_ VGND VGND VPWR VPWR _2530_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4300_ _3127_ _3402_ _3405_ _1701_ VGND VGND VPWR VPWR _3406_ sky130_fd_sc_hd__o211a_1
X_5280_ _0583_ _0584_ _1734_ _3580_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__a31o_1
XFILLER_0_51_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4231_ _3262_ _3336_ VGND VGND VPWR VPWR _3338_ sky130_fd_sc_hd__or2_1
X_4162_ _3269_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_2
X_4093_ _0063_ _3161_ VGND VGND VPWR VPWR _3201_ sky130_fd_sc_hd__and2_2
XFILLER_0_148_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4995_ _0392_ _0393_ _0371_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__a21oi_1
X_6803_ _2180_ _2181_ VGND VGND VPWR VPWR _2371_ sky130_fd_sc_hd__or2b_1
XFILLER_0_148_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3946_ _1023_ _2346_ _2029_ VGND VGND VPWR VPWR _2357_ sky130_fd_sc_hd__mux2_2
XFILLER_0_58_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6734_ _1953_ _1960_ _2295_ VGND VGND VPWR VPWR _2296_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_555 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3877_ _0881_ _0521_ _1056_ _1002_ VGND VGND VPWR VPWR _1603_ sky130_fd_sc_hd__and4_1
XFILLER_0_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6665_ _2664_ _0327_ _0454_ _2259_ VGND VGND VPWR VPWR _2220_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_131_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6596_ _1745_ _2142_ _2143_ VGND VGND VPWR VPWR _2144_ sky130_fd_sc_hd__a21bo_1
X_5616_ _3644_ _0339_ _0340_ _2434_ VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5547_ _0824_ _0895_ _0997_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__o21ai_1
X_5478_ _0919_ _0920_ _0898_ _0899_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__o211a_1
X_4429_ _3531_ _2368_ _2423_ _0161_ VGND VGND VPWR VPWR _3533_ sky130_fd_sc_hd__a22o_1
X_7217_ _2581_ _2582_ VGND VGND VPWR VPWR _2824_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7148_ _2746_ _2747_ VGND VGND VPWR VPWR _2748_ sky130_fd_sc_hd__xnor2_1
X_7079_ _2301_ _2306_ _2300_ VGND VGND VPWR VPWR _2673_ sky130_fd_sc_hd__a21o_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_773 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4780_ _0092_ _0159_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__xnor2_2
X_3800_ _0368_ _0728_ _0750_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__o21a_1
XFILLER_0_68_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6450_ _1982_ _1983_ VGND VGND VPWR VPWR _1984_ sky130_fd_sc_hd__and2_1
XFILLER_0_140_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5401_ _3582_ _3584_ _0199_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__mux2_1
X_6381_ _1735_ net201 _1907_ _1908_ VGND VGND VPWR VPWR _1910_ sky130_fd_sc_hd__o211a_4
XFILLER_0_30_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5332_ _0754_ _0762_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5263_ _0654_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__clkbuf_4
X_4214_ _3241_ _3244_ _3243_ VGND VGND VPWR VPWR _3321_ sky130_fd_sc_hd__a21bo_1
X_5194_ _0609_ _0610_ _0480_ _0482_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7002_ _2675_ _2718_ _0328_ _0559_ _2426_ VGND VGND VPWR VPWR _2589_ sky130_fd_sc_hd__a41o_1
X_4145_ _3250_ _3251_ _3252_ VGND VGND VPWR VPWR _3253_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4076_ _3174_ _3184_ VGND VGND VPWR VPWR _3185_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_92_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4978_ _2653_ _0374_ _0375_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6717_ _2126_ net177 _2275_ _2276_ _3192_ VGND VGND VPWR VPWR _2277_ sky130_fd_sc_hd__a311o_1
XFILLER_0_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3929_ _2160_ VGND VGND VPWR VPWR _2171_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_117_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6648_ _0117_ net48 _2198_ _2199_ VGND VGND VPWR VPWR _2201_ sky130_fd_sc_hd__nand4_2
XFILLER_0_33_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6579_ _2125_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_6
XFILLER_0_100_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_731 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_810 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5950_ net133 _1138_ _1139_ VGND VGND VPWR VPWR _1438_ sky130_fd_sc_hd__nand3_1
XFILLER_0_153_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4901_ _0220_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5881_ _1224_ _1218_ VGND VGND VPWR VPWR _1363_ sky130_fd_sc_hd__and2b_1
XFILLER_0_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4832_ _0739_ _0423_ _3718_ _0099_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__and4_1
XFILLER_0_8_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4763_ _0048_ _0049_ _0050_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4694_ _0029_ _0065_ _0066_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__or3_4
X_7482_ _0860_ _0850_ _3107_ _0368_ _3109_ VGND VGND VPWR VPWR _3110_ sky130_fd_sc_hd__o221a_1
X_6502_ _1895_ _1897_ _1894_ VGND VGND VPWR VPWR _2042_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_15_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6433_ _1676_ _1792_ _1811_ VGND VGND VPWR VPWR _1966_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_141_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6364_ _2259_ _0220_ _1889_ _1890_ VGND VGND VPWR VPWR _1891_ sky130_fd_sc_hd__nand4_1
XFILLER_0_3_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5315_ _0611_ _0612_ _0646_ _0647_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__or4_4
X_6295_ _1672_ _1674_ VGND VGND VPWR VPWR _1815_ sky130_fd_sc_hd__and2_1
X_5246_ _0667_ _0668_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5177_ _0490_ _0500_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__nand2_1
X_4128_ _3169_ _1264_ _0314_ _0030_ VGND VGND VPWR VPWR _3236_ sky130_fd_sc_hd__a22oi_2
X_4059_ _1449_ _1493_ VGND VGND VPWR VPWR _3168_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_751 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5100_ _3451_ _3452_ _0380_ _2489_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__nand4_1
X_6080_ _1541_ _1542_ _1577_ _1578_ VGND VGND VPWR VPWR _1580_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_0_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5031_ _3702_ _0433_ _0429_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__mux2_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6982_ _2431_ VGND VGND VPWR VPWR _2567_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5933_ _1381_ _1382_ _1418_ _1419_ VGND VGND VPWR VPWR _1420_ sky130_fd_sc_hd__nor4_2
XFILLER_0_146_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5864_ _1342_ _1343_ _2313_ net41 VGND VGND VPWR VPWR _1344_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_8_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4815_ _3486_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5795_ _1151_ _1267_ _1155_ _3192_ VGND VGND VPWR VPWR _1269_ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4746_ _0043_ _0044_ _0045_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_16_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4677_ _0281_ _3537_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__and2_1
X_7465_ _0259_ _0576_ VGND VGND VPWR VPWR _3092_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7396_ _2949_ _3018_ VGND VGND VPWR VPWR _3019_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6416_ _3571_ _1937_ _1938_ _1947_ VGND VGND VPWR VPWR _1948_ sky130_fd_sc_hd__a31o_1
X_6347_ _1725_ _1727_ VGND VGND VPWR VPWR _1872_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6278_ _1648_ _1649_ _1645_ VGND VGND VPWR VPWR _1796_ sky130_fd_sc_hd__o21ai_1
X_5229_ _0524_ _0526_ net113 _0649_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_79_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_838 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4600_ _3283_ _3702_ _3087_ VGND VGND VPWR VPWR _3703_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5580_ _0919_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4531_ _2302_ _3632_ _3633_ _0085_ VGND VGND VPWR VPWR _3634_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4462_ _3476_ _3564_ _3565_ VGND VGND VPWR VPWR _3566_ sky130_fd_sc_hd__and3_1
X_7250_ _2660_ _2859_ VGND VGND VPWR VPWR _2860_ sky130_fd_sc_hd__nand2_1
X_6201_ _1887_ _1710_ _1711_ VGND VGND VPWR VPWR _1713_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4393_ _3482_ _3497_ _3265_ VGND VGND VPWR VPWR _3498_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7181_ _2782_ _2783_ VGND VGND VPWR VPWR _2785_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6132_ _1634_ _1636_ VGND VGND VPWR VPWR _1637_ sky130_fd_sc_hd__nor2_1
X_6063_ _1558_ _1560_ _1561_ VGND VGND VPWR VPWR _1562_ sky130_fd_sc_hd__nand3_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ _0207_ _0285_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6965_ _3513_ _2609_ _1865_ _3424_ VGND VGND VPWR VPWR _2548_ sky130_fd_sc_hd__a22o_1
X_5916_ _0488_ _0390_ _1887_ net15 VGND VGND VPWR VPWR _1401_ sky130_fd_sc_hd__nand4_1
XFILLER_0_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6896_ _2448_ _2449_ _2471_ _2472_ VGND VGND VPWR VPWR _2473_ sky130_fd_sc_hd__nor4_1
XFILLER_0_36_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5847_ _0434_ net46 _1294_ _0466_ VGND VGND VPWR VPWR _1325_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5778_ _1247_ _1248_ _1119_ _1121_ VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4729_ net64 VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_72_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7448_ _3587_ _3073_ VGND VGND VPWR VPWR _3074_ sky130_fd_sc_hd__nand2_2
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7379_ _2994_ _2999_ VGND VGND VPWR VPWR _3000_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6750_ _2007_ _1821_ _1810_ _1778_ _0583_ _0584_ VGND VGND VPWR VPWR _2312_ sky130_fd_sc_hd__mux4_1
XFILLER_0_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3962_ _2521_ VGND VGND VPWR VPWR _2532_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5701_ _1163_ _1164_ VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3893_ _1767_ VGND VGND VPWR VPWR _1778_ sky130_fd_sc_hd__buf_4
XFILLER_0_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6681_ _2235_ _2236_ VGND VGND VPWR VPWR _2238_ sky130_fd_sc_hd__or2b_1
XFILLER_0_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5632_ _0956_ _0975_ _0976_ VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__nand3_2
XFILLER_0_72_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5563_ _1011_ _1014_ VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4514_ _0314_ net64 _3572_ net163 VGND VGND VPWR VPWR _3617_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7302_ _2913_ _2915_ VGND VGND VPWR VPWR _2916_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5494_ _0938_ _0939_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_41_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4445_ _3545_ _3546_ _3547_ VGND VGND VPWR VPWR _3549_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7233_ _2838_ _2840_ _2638_ _2640_ VGND VGND VPWR VPWR _2842_ sky130_fd_sc_hd__a211oi_2
X_4376_ _2171_ _3425_ VGND VGND VPWR VPWR _3481_ sky130_fd_sc_hd__nor2_1
X_7164_ _2763_ _2764_ _2705_ _2706_ VGND VGND VPWR VPWR _2766_ sky130_fd_sc_hd__a211o_1
XFILLER_0_1_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6115_ _1437_ _1441_ _1597_ VGND VGND VPWR VPWR _1618_ sky130_fd_sc_hd__or3_4
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7095_ _2682_ _2685_ _2690_ VGND VGND VPWR VPWR _2691_ sky130_fd_sc_hd__or3_1
X_6046_ _1394_ _1413_ _1414_ VGND VGND VPWR VPWR _1543_ sky130_fd_sc_hd__nor3_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6948_ _3386_ _1898_ VGND VGND VPWR VPWR _2529_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6879_ _2244_ _2253_ VGND VGND VPWR VPWR _2454_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4230_ _3262_ _3336_ VGND VGND VPWR VPWR _3337_ sky130_fd_sc_hd__nand2_1
X_4161_ _3206_ _3230_ _3268_ VGND VGND VPWR VPWR _3269_ sky130_fd_sc_hd__or3_1
X_4092_ _0980_ _0969_ _0870_ VGND VGND VPWR VPWR _3200_ sky130_fd_sc_hd__o21a_2
XFILLER_0_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6802_ _2366_ _2367_ _2151_ _2334_ VGND VGND VPWR VPWR _2370_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_148_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4994_ _0371_ _0392_ _0393_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6733_ _1949_ _1810_ VGND VGND VPWR VPWR _2295_ sky130_fd_sc_hd__and2b_1
X_3945_ _2335_ VGND VGND VPWR VPWR _2346_ sky130_fd_sc_hd__buf_6
XFILLER_0_147_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6664_ _2259_ _2653_ _0326_ _0453_ VGND VGND VPWR VPWR _2219_ sky130_fd_sc_hd__and4_1
X_5615_ _0948_ _0955_ VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__and2_1
X_3876_ _1012_ _1581_ VGND VGND VPWR VPWR _1592_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6595_ _0052_ net16 net17 _0172_ VGND VGND VPWR VPWR _2143_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5546_ _0995_ _0996_ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5477_ _0898_ _0899_ _0919_ _0920_ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4428_ _0161_ _3531_ _2368_ VGND VGND VPWR VPWR _3532_ sky130_fd_sc_hd__and3_1
X_7216_ _2628_ _2636_ VGND VGND VPWR VPWR _2823_ sky130_fd_sc_hd__nand2_1
X_4359_ _3439_ _3462_ _3463_ VGND VGND VPWR VPWR _3464_ sky130_fd_sc_hd__nand3_4
X_7147_ _0293_ _2510_ VGND VGND VPWR VPWR _2747_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7078_ _2670_ _2671_ VGND VGND VPWR VPWR _2672_ sky130_fd_sc_hd__nor2_2
X_6029_ _2259_ _3718_ _0099_ _2204_ VGND VGND VPWR VPWR _1524_ sky130_fd_sc_hd__a22o_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6380_ _1884_ _1885_ _1905_ _1906_ VGND VGND VPWR VPWR _1908_ sky130_fd_sc_hd__o22ai_4
X_5400_ _0829_ _0834_ _0835_ _0836_ _3596_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__a311o_1
XFILLER_0_140_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5331_ _0759_ _0760_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5262_ _0592_ _0557_ _0684_ _3192_ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__a31o_1
X_7001_ _2421_ _2429_ VGND VGND VPWR VPWR _2588_ sky130_fd_sc_hd__nand2_1
X_4213_ _3317_ _3318_ _3316_ VGND VGND VPWR VPWR _3320_ sky130_fd_sc_hd__a21o_1
X_5193_ _0480_ _0482_ _0609_ _0610_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_76_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4144_ _3174_ _3183_ _3182_ VGND VGND VPWR VPWR _3252_ sky130_fd_sc_hd__o21bai_4
X_4075_ _3182_ _3183_ VGND VGND VPWR VPWR _3184_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4977_ net191 net3 _2642_ _3169_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__a22o_1
X_6716_ _2126_ net177 _2275_ VGND VGND VPWR VPWR _2276_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3928_ _2149_ VGND VGND VPWR VPWR _2160_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3859_ _0183_ _1384_ _1395_ VGND VGND VPWR VPWR _1406_ sky130_fd_sc_hd__nand3_1
XFILLER_0_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6647_ _0117_ net48 _2198_ _2199_ VGND VGND VPWR VPWR _2200_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_468 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6578_ _2113_ _2118_ _2124_ VGND VGND VPWR VPWR _2125_ sky130_fd_sc_hd__or3b_4
X_5529_ _0975_ _0976_ _0956_ VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_30_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4900_ _0287_ _0289_ _3192_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5880_ _1202_ _1211_ VGND VGND VPWR VPWR _1361_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_527 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4831_ _0335_ _3718_ _0100_ _0423_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4762_ _0137_ _0138_ _0136_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4693_ _0062_ _0064_ _3662_ _0031_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__o211a_1
X_7481_ _0270_ net123 _1187_ _0368_ VGND VGND VPWR VPWR _3109_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_71_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6501_ _3620_ _2784_ _2037_ _2038_ VGND VGND VPWR VPWR _2041_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_125_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6432_ _1918_ VGND VGND VPWR VPWR _1965_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6363_ _3718_ _2696_ _0100_ _2653_ VGND VGND VPWR VPWR _1890_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5314_ _0646_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6294_ _1678_ _1680_ _1739_ _1740_ VGND VGND VPWR VPWR _1814_ sky130_fd_sc_hd__nor4_1
X_5245_ _0484_ _0486_ _0666_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5176_ _0540_ _0541_ _0542_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__nand3_1
X_4127_ _3233_ _3234_ VGND VGND VPWR VPWR _3235_ sky130_fd_sc_hd__or2_4
XFILLER_0_127_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4058_ _2980_ _3002_ _3013_ _3166_ VGND VGND VPWR VPWR _3167_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _3135_ _3134_ _3133_ _2675_ _3046_ _3591_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__mux4_2
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6981_ _2562_ _2563_ _2369_ _2395_ VGND VGND VPWR VPWR _2566_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_88_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5932_ _1415_ _1416_ _1245_ _1383_ VGND VGND VPWR VPWR _1419_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_76_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5863_ _2434_ _0325_ _0452_ _3442_ VGND VGND VPWR VPWR _1343_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_8_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5794_ _1151_ _1155_ _1267_ VGND VGND VPWR VPWR _1268_ sky130_fd_sc_hd__a21oi_1
X_4814_ _3194_ _0191_ _0192_ _3414_ _0197_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4745_ _0106_ _3386_ _0036_ _0035_ _2324_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__a32o_1
XFILLER_0_56_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4676_ _0043_ _0046_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7464_ _0259_ _0576_ VGND VGND VPWR VPWR _3091_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7395_ _2992_ _3017_ VGND VGND VPWR VPWR _3018_ sky130_fd_sc_hd__xnor2_1
X_6415_ _1766_ _1943_ _1944_ _1946_ VGND VGND VPWR VPWR _1947_ sky130_fd_sc_hd__or4b_1
XFILLER_0_102_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6346_ _1867_ _1868_ _1869_ VGND VGND VPWR VPWR _1871_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6277_ _1650_ _1658_ VGND VGND VPWR VPWR _1795_ sky130_fd_sc_hd__or2_1
X_5228_ _0611_ _0612_ _0646_ _0647_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__o22a_1
X_5159_ _0571_ _0572_ _0573_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_560 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4530_ _3270_ VGND VGND VPWR VPWR _3633_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4461_ _3563_ _3561_ _3562_ VGND VGND VPWR VPWR _3565_ sky130_fd_sc_hd__nand3_1
XFILLER_0_13_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6200_ _0030_ net13 net14 _3169_ VGND VGND VPWR VPWR _1711_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7180_ _2774_ _2781_ VGND VGND VPWR VPWR _2783_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4392_ _3389_ _3391_ _3496_ VGND VGND VPWR VPWR _3497_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6131_ _1629_ _1630_ _1633_ VGND VGND VPWR VPWR _1636_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _1402_ _1403_ _1401_ VGND VGND VPWR VPWR _1561_ sky130_fd_sc_hd__a21bo_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _0321_ _0414_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6964_ _2545_ _2546_ VGND VGND VPWR VPWR _2547_ sky130_fd_sc_hd__xor2_2
X_5915_ _1398_ _1399_ VGND VGND VPWR VPWR _1400_ sky130_fd_sc_hd__xor2_1
X_6895_ _2469_ _2470_ _2451_ _2452_ VGND VGND VPWR VPWR _2472_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5846_ _1191_ _1192_ _1254_ net204 VGND VGND VPWR VPWR _1324_ sky130_fd_sc_hd__nor4_2
XFILLER_0_8_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5777_ _1119_ net128 _1247_ _1248_ VGND VGND VPWR VPWR _1249_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_16_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4728_ _0101_ _0102_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4659_ _0018_ _0027_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__xnor2_1
X_7447_ _3400_ _3403_ _3072_ _3401_ _0861_ _0867_ VGND VGND VPWR VPWR _3073_ sky130_fd_sc_hd__mux4_1
XFILLER_0_142_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7378_ _2995_ _2998_ VGND VGND VPWR VPWR _2999_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6329_ _3451_ _3452_ net17 net18 VGND VGND VPWR VPWR _1852_ sky130_fd_sc_hd__nand4_2
XFILLER_0_87_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_530 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3961_ net9 VGND VGND VPWR VPWR _2521_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_147_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5700_ _0707_ _1007_ _1161_ _1162_ VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__a22oi_1
X_3892_ net18 VGND VGND VPWR VPWR _1767_ sky130_fd_sc_hd__buf_2
X_6680_ _2191_ _2192_ _2233_ _2234_ VGND VGND VPWR VPWR _2236_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_727 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5631_ _1086_ _1087_ _1070_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5562_ _0878_ _1001_ _1013_ VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__a21o_1
X_4513_ _0314_ _0412_ net64 _3572_ VGND VGND VPWR VPWR _3616_ sky130_fd_sc_hd__and4_1
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7301_ _3139_ _1608_ _2802_ net102 VGND VGND VPWR VPWR _2915_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_41_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5493_ _0755_ _0756_ _0757_ VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_14_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7232_ _2638_ _2640_ _2838_ _2840_ VGND VGND VPWR VPWR _2841_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4444_ _3545_ _3546_ _3547_ VGND VGND VPWR VPWR _3548_ sky130_fd_sc_hd__nand3_2
XFILLER_0_1_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7163_ _2705_ _2706_ _2763_ _2764_ VGND VGND VPWR VPWR _2765_ sky130_fd_sc_hd__o211ai_4
X_4375_ _2171_ _3425_ VGND VGND VPWR VPWR _3480_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7094_ _3156_ _0201_ _2689_ _0844_ VGND VGND VPWR VPWR _2690_ sky130_fd_sc_hd__a2bb2o_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6114_ _0419_ _1615_ _1616_ VGND VGND VPWR VPWR _1617_ sky130_fd_sc_hd__and3_1
X_6045_ _1539_ _1540_ _1520_ _1521_ VGND VGND VPWR VPWR _1542_ sky130_fd_sc_hd__o211a_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6947_ _2526_ _2527_ VGND VGND VPWR VPWR _2528_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6878_ _2252_ _2245_ VGND VGND VPWR VPWR _2453_ sky130_fd_sc_hd__or2b_1
XFILLER_0_37_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5829_ _1011_ _1027_ _1272_ _1304_ _1271_ VGND VGND VPWR VPWR _1305_ sky130_fd_sc_hd__o311ai_4
XFILLER_0_9_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_474 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4160_ _1668_ _3261_ _3262_ _3267_ VGND VGND VPWR VPWR _3268_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4091_ _2412_ _3198_ VGND VGND VPWR VPWR _3199_ sky130_fd_sc_hd__and2_1
X_6801_ _2151_ _2334_ _2366_ _2367_ VGND VGND VPWR VPWR _2369_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4993_ _0388_ _0389_ _0391_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3944_ _2324_ VGND VGND VPWR VPWR _2335_ sky130_fd_sc_hd__buf_4
XFILLER_0_19_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6732_ _3156_ _3699_ _2288_ _2290_ _2293_ VGND VGND VPWR VPWR _2294_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3875_ _1351_ _1340_ VGND VGND VPWR VPWR _1581_ sky130_fd_sc_hd__and2b_1
X_6663_ _2032_ _2035_ _2033_ VGND VGND VPWR VPWR _2218_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_45_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5614_ _0954_ _0949_ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__and2b_1
XFILLER_0_61_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6594_ _0172_ _0052_ net16 VGND VGND VPWR VPWR _2142_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5545_ net140 _0815_ _0814_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__a21o_1
X_5476_ _0764_ _0900_ _0918_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4427_ net59 VGND VGND VPWR VPWR _3531_ sky130_fd_sc_hd__clkbuf_4
X_7215_ _2635_ _2629_ VGND VGND VPWR VPWR _2822_ sky130_fd_sc_hd__or2b_1
XFILLER_0_111_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7146_ _2744_ _2745_ VGND VGND VPWR VPWR _2746_ sky130_fd_sc_hd__or2_1
X_4358_ _3459_ _3460_ _3461_ VGND VGND VPWR VPWR _3463_ sky130_fd_sc_hd__a21o_1
X_4289_ _3274_ _3394_ VGND VGND VPWR VPWR _3395_ sky130_fd_sc_hd__nor2_1
X_7077_ _2018_ net54 VGND VGND VPWR VPWR _2671_ sky130_fd_sc_hd__nor2_1
X_6028_ _2215_ _2259_ _0099_ VGND VGND VPWR VPWR _1523_ sky130_fd_sc_hd__and3_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5330_ _0601_ _0602_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5261_ _0592_ _0557_ _0684_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4212_ _3316_ _3317_ _3318_ VGND VGND VPWR VPWR _3319_ sky130_fd_sc_hd__nand3_1
X_7000_ _2584_ _2585_ VGND VGND VPWR VPWR _2586_ sky130_fd_sc_hd__and2_1
X_5192_ _0497_ _0593_ _0607_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__and3_1
X_4143_ _3248_ _3249_ _3240_ VGND VGND VPWR VPWR _3251_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4074_ _3179_ _3180_ _3181_ VGND VGND VPWR VPWR _3183_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_558 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4976_ _3352_ _0373_ net3 VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__and3_1
X_6715_ _2102_ _2274_ VGND VGND VPWR VPWR _2275_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3927_ net32 VGND VGND VPWR VPWR _2149_ sky130_fd_sc_hd__buf_4
XFILLER_0_73_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3858_ _1329_ _1362_ VGND VGND VPWR VPWR _1395_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6646_ _2324_ _2390_ _1169_ _1294_ VGND VGND VPWR VPWR _2199_ sky130_fd_sc_hd__nand4_2
XFILLER_0_46_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3789_ net66 net67 net68 VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__or3_4
XFILLER_0_15_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6577_ _3156_ _3585_ _2123_ VGND VGND VPWR VPWR _2124_ sky130_fd_sc_hd__o21a_1
XFILLER_0_132_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5528_ _0956_ _0975_ _0976_ VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5459_ _1056_ _0722_ _0875_ _1002_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__a22o_1
X_7129_ _3386_ _1898_ _2528_ _2527_ VGND VGND VPWR VPWR _2727_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4830_ _0122_ _0129_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4761_ _0136_ _0137_ _0138_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__nand3_1
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4692_ _3662_ _0031_ _0062_ _0064_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__a211oi_2
X_7480_ _0750_ _3158_ _3204_ VGND VGND VPWR VPWR _3107_ sky130_fd_sc_hd__a21oi_1
X_6500_ _3620_ _2784_ _2037_ _2038_ VGND VGND VPWR VPWR _2039_ sky130_fd_sc_hd__and4_1
XFILLER_0_7_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6431_ _1923_ _1924_ VGND VGND VPWR VPWR _1964_ sky130_fd_sc_hd__nor2_2
XFILLER_0_140_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6362_ _2707_ _0100_ _3722_ VGND VGND VPWR VPWR _1889_ sky130_fd_sc_hd__nand3_1
XFILLER_0_140_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5313_ _0458_ _0662_ _0738_ _0740_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__nand4_2
XFILLER_0_87_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6293_ _1791_ _1812_ VGND VGND VPWR VPWR _1813_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5244_ _0484_ _0486_ _0666_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__o21ai_1
X_5175_ _0320_ _0556_ _0557_ _0591_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__a31o_2
X_4126_ _0466_ _3197_ _3171_ _3232_ VGND VGND VPWR VPWR _3234_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_39_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4057_ _0838_ _3097_ _3126_ _3157_ _3165_ VGND VGND VPWR VPWR _3166_ sky130_fd_sc_hd__a311o_1
XFILLER_0_78_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4959_ _0334_ _0336_ _0353_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__nor3_1
XFILLER_0_47_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6629_ _2178_ _2179_ VGND VGND VPWR VPWR _2180_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_552 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_815 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6980_ _2369_ _2395_ _2562_ _2563_ VGND VGND VPWR VPWR _2564_ sky130_fd_sc_hd__o211a_1
X_5931_ _1245_ _1383_ _1415_ _1416_ VGND VGND VPWR VPWR _1418_ sky130_fd_sc_hd__o211a_4
XFILLER_0_76_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5862_ _2368_ _2423_ _0325_ _0452_ VGND VGND VPWR VPWR _1342_ sky130_fd_sc_hd__and4_1
XFILLER_0_146_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5793_ _1265_ _1266_ VGND VGND VPWR VPWR _1267_ sky130_fd_sc_hd__xor2_2
XFILLER_0_75_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4813_ _0176_ _0193_ _0196_ _3201_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4744_ _0040_ _0060_ _0061_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__nand3_2
XFILLER_0_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4675_ _0044_ _0045_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7463_ _0237_ _0309_ _3712_ _0248_ _3089_ VGND VGND VPWR VPWR _3090_ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7394_ _3000_ _3016_ VGND VGND VPWR VPWR _3017_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6414_ _3156_ _3493_ _1928_ _1945_ VGND VGND VPWR VPWR _1946_ sky130_fd_sc_hd__o22a_1
XFILLER_0_43_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6345_ _1867_ _1868_ _1869_ VGND VGND VPWR VPWR _1870_ sky130_fd_sc_hd__and3_4
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6276_ _1655_ _1656_ VGND VGND VPWR VPWR _1794_ sky130_fd_sc_hd__nand2_1
X_5227_ _0611_ _0612_ _0646_ _0647_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__nor4_1
X_5158_ _0838_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__clkbuf_4
X_4109_ _3215_ _3216_ VGND VGND VPWR VPWR _3217_ sky130_fd_sc_hd__xnor2_1
X_5089_ _0492_ _0495_ _0496_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__or3_4
XFILLER_0_98_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_699 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4460_ _3561_ _3562_ _3563_ VGND VGND VPWR VPWR _3564_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_636 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4391_ _3386_ _2138_ VGND VGND VPWR VPWR _3496_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6130_ _1629_ _1630_ _1633_ VGND VGND VPWR VPWR _1634_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _1555_ _1556_ _1557_ VGND VGND VPWR VPWR _1560_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _0410_ _0413_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__xnor2_2
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6963_ _0293_ _2784_ VGND VGND VPWR VPWR _2546_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5914_ _0042_ _2532_ VGND VGND VPWR VPWR _1399_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6894_ _2451_ _2452_ _2469_ _2470_ VGND VGND VPWR VPWR _2471_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5845_ _1320_ _1322_ VGND VGND VPWR VPWR _1323_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5776_ _1245_ _1246_ _1226_ VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_8_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4727_ _0707_ _0466_ _3719_ _0100_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__and4_1
X_4658_ _0019_ _0026_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__xnor2_1
X_7446_ _2357_ _3070_ _2467_ _3071_ _0866_ _0864_ VGND VGND VPWR VPWR _3072_ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4589_ _3688_ _3690_ VGND VGND VPWR VPWR _3692_ sky130_fd_sc_hd__and2_1
X_7377_ _2996_ _2997_ VGND VGND VPWR VPWR _2998_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6328_ _1720_ _1721_ _1731_ VGND VGND VPWR VPWR _1851_ sky130_fd_sc_hd__nor3_2
XFILLER_0_110_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6259_ _0878_ _1775_ _1013_ VGND VGND VPWR VPWR _1776_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3960_ _2499_ VGND VGND VPWR VPWR _2510_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3891_ _1745_ VGND VGND VPWR VPWR _1756_ sky130_fd_sc_hd__buf_4
XFILLER_0_73_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5630_ _1070_ _1086_ _1087_ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__nor3_1
XFILLER_0_116_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5561_ _0875_ _0862_ VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__and2b_1
XFILLER_0_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4512_ _3522_ _3527_ _3614_ VGND VGND VPWR VPWR _3615_ sky130_fd_sc_hd__o21ai_2
X_5492_ _0935_ _0937_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7300_ _2802_ net102 _3139_ _1608_ VGND VGND VPWR VPWR _2913_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7231_ _2836_ _2837_ _2822_ _2823_ VGND VGND VPWR VPWR _2840_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_123_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4443_ _3446_ _3458_ _3457_ VGND VGND VPWR VPWR _3547_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_110_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4374_ _3384_ _3475_ VGND VGND VPWR VPWR _3479_ sky130_fd_sc_hd__or2_4
XFILLER_0_95_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7162_ _2739_ _2741_ _2760_ _2761_ VGND VGND VPWR VPWR _2764_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7093_ _3097_ _0188_ _1284_ _2688_ _0867_ _0573_ VGND VGND VPWR VPWR _2689_ sky130_fd_sc_hd__mux4_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6113_ _1611_ _1614_ VGND VGND VPWR VPWR _1616_ sky130_fd_sc_hd__or2_1
X_6044_ _1520_ _1521_ _1539_ _1540_ VGND VGND VPWR VPWR _1541_ sky130_fd_sc_hd__a211oi_4
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6946_ _3197_ _3273_ _1931_ _1952_ VGND VGND VPWR VPWR _2527_ sky130_fd_sc_hd__and4_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6877_ _2255_ _2257_ VGND VGND VPWR VPWR _2452_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5828_ _1010_ _1270_ VGND VGND VPWR VPWR _1304_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5759_ _2565_ _1227_ _1228_ VGND VGND VPWR VPWR _1229_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_9_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_444 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7429_ _0717_ net123 _1187_ _0685_ _3053_ VGND VGND VPWR VPWR _3054_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4090_ _3197_ VGND VGND VPWR VPWR _3198_ sky130_fd_sc_hd__buf_2
XFILLER_0_65_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6800_ _2353_ _2354_ _2365_ VGND VGND VPWR VPWR _2367_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_147_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4992_ _0388_ _0389_ _0391_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__nand3_2
XFILLER_0_147_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3943_ _2313_ VGND VGND VPWR VPWR _2324_ sky130_fd_sc_hd__buf_4
X_6731_ _2121_ _2291_ VGND VGND VPWR VPWR _2293_ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3874_ _1548_ _1559_ VGND VGND VPWR VPWR _1570_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6662_ _2075_ _2077_ VGND VGND VPWR VPWR _2217_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5613_ _0935_ _0937_ _0939_ _1069_ VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__o31a_1
XFILLER_0_61_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6593_ _2136_ _2137_ _2139_ VGND VGND VPWR VPWR _2141_ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5544_ _0993_ _0994_ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__or2b_4
XFILLER_0_14_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5475_ _0764_ _0900_ _0918_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_14_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4426_ _2423_ VGND VGND VPWR VPWR _3530_ sky130_fd_sc_hd__buf_4
XFILLER_0_69_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7214_ _2819_ _2820_ VGND VGND VPWR VPWR _2821_ sky130_fd_sc_hd__nand2_1
X_7145_ _3720_ _0174_ _2543_ _2576_ VGND VGND VPWR VPWR _2745_ sky130_fd_sc_hd__and4_1
X_4357_ _3459_ _3460_ _3461_ VGND VGND VPWR VPWR _3462_ sky130_fd_sc_hd__nand3_4
X_4288_ _2456_ _3273_ _2401_ _3198_ VGND VGND VPWR VPWR _3394_ sky130_fd_sc_hd__o211a_1
X_7076_ _2018_ net54 VGND VGND VPWR VPWR _2670_ sky130_fd_sc_hd__and2_2
X_6027_ _1385_ _1392_ _1391_ VGND VGND VPWR VPWR _1522_ sky130_fd_sc_hd__a21o_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6929_ _2504_ _2505_ _2506_ VGND VGND VPWR VPWR _2508_ sky130_fd_sc_hd__nand3_1
XFILLER_0_77_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5260_ _0681_ _0683_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4211_ net44 net29 net30 net33 VGND VGND VPWR VPWR _3318_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5191_ _0497_ _0593_ _0607_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__a21oi_4
X_4142_ _3240_ _3248_ _3249_ VGND VGND VPWR VPWR _3250_ sky130_fd_sc_hd__nand3_1
X_4073_ _3179_ _3180_ _3181_ VGND VGND VPWR VPWR _3182_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4975_ net59 VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3926_ _2127_ VGND VGND VPWR VPWR _2138_ sky130_fd_sc_hd__clkbuf_4
X_6714_ _2128_ _2273_ VGND VGND VPWR VPWR _2274_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_73_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3857_ _1002_ VGND VGND VPWR VPWR _1384_ sky130_fd_sc_hd__buf_4
XFILLER_0_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6645_ _2390_ _1169_ _1294_ _2324_ VGND VGND VPWR VPWR _2198_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3788_ net65 VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6576_ _1950_ _2120_ _2122_ VGND VGND VPWR VPWR _2123_ sky130_fd_sc_hd__o21ba_1
X_5527_ _0972_ _0973_ _0974_ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5458_ _0745_ _0746_ _0764_ _0765_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_2_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5389_ _3192_ _0824_ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__or2_1
X_4409_ _3512_ VGND VGND VPWR VPWR _3513_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7128_ _2722_ _2723_ _2724_ VGND VGND VPWR VPWR _2726_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7059_ _2610_ _2611_ _2649_ _2650_ VGND VGND VPWR VPWR _2651_ sky130_fd_sc_hd__nand4_2
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_695 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4760_ _3449_ _3448_ _2642_ _2686_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__nand4_2
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4691_ _0060_ _0061_ _0040_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6430_ _1953_ _1960_ _1961_ VGND VGND VPWR VPWR _1962_ sky130_fd_sc_hd__o21a_1
XFILLER_0_102_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6361_ _1722_ _1730_ VGND VGND VPWR VPWR _1888_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5312_ _0458_ _0662_ _0738_ _0740_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6292_ _1793_ _1811_ VGND VGND VPWR VPWR _1812_ sky130_fd_sc_hd__xnor2_1
X_5243_ _0662_ _0665_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__xnor2_1
X_5174_ _3571_ _0568_ _0577_ _0590_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__a211o_1
X_4125_ _3171_ _3232_ net1 _3197_ VGND VGND VPWR VPWR _3233_ sky130_fd_sc_hd__o211a_1
X_4056_ _1187_ _2914_ _2925_ _1176_ _3164_ VGND VGND VPWR VPWR _3165_ sky130_fd_sc_hd__a221o_1
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4958_ _0334_ _0336_ _0353_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__o21a_1
X_4889_ _0277_ _0278_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__nor2_2
X_3909_ net16 VGND VGND VPWR VPWR _1952_ sky130_fd_sc_hd__buf_2
XFILLER_0_61_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6628_ _3620_ _2510_ VGND VGND VPWR VPWR _2179_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6559_ _2102_ _2103_ VGND VGND VPWR VPWR _2104_ sky130_fd_sc_hd__and2_2
XFILLER_0_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_776 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5930_ _1413_ _1414_ _1394_ VGND VGND VPWR VPWR _1416_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5861_ _1175_ _1178_ VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5792_ net132 _1139_ _1138_ VGND VGND VPWR VPWR _1266_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_91_808 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4812_ _0195_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__buf_2
XFILLER_0_8_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4743_ _0116_ _0118_ _0094_ _0096_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7462_ _0860_ _0869_ _3088_ _0674_ VGND VGND VPWR VPWR _3089_ sky130_fd_sc_hd__o22a_1
XFILLER_0_71_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4674_ _0161_ _3531_ _2106_ net32 VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__and4_1
X_6413_ _3589_ _1929_ _0000_ VGND VGND VPWR VPWR _1945_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_43_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_779 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7393_ _3006_ _3015_ VGND VGND VPWR VPWR _3016_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_141_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6344_ _1709_ _1715_ _1708_ VGND VGND VPWR VPWR _1869_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6275_ _1676_ _1792_ VGND VGND VPWR VPWR _1793_ sky130_fd_sc_hd__nand2_1
X_5226_ _0644_ _0645_ _0519_ _0613_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5157_ _3401_ _3403_ _0199_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__mux2_1
X_4108_ _3159_ _2991_ _2914_ VGND VGND VPWR VPWR _3216_ sky130_fd_sc_hd__a21oi_1
X_5088_ _0493_ _0494_ _3388_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__a21oi_1
X_4039_ _3146_ _3147_ _0947_ VGND VGND VPWR VPWR _3148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_746 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4390_ _3127_ _3491_ _3494_ _1701_ VGND VGND VPWR VPWR _3495_ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _1555_ _1556_ _1557_ VGND VGND VPWR VPWR _1558_ sky130_fd_sc_hd__nand3_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _0283_ _0282_ _0411_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__o21ai_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6962_ _2543_ _2542_ _2544_ VGND VGND VPWR VPWR _2545_ sky130_fd_sc_hd__a21bo_1
X_5913_ _2598_ _1396_ _1397_ VGND VGND VPWR VPWR _1398_ sky130_fd_sc_hd__a21bo_1
X_6893_ _2466_ _2468_ _2453_ _2454_ VGND VGND VPWR VPWR _2470_ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5844_ _3209_ _1170_ _1168_ _1321_ VGND VGND VPWR VPWR _1322_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_8_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5775_ _1226_ _1245_ _1246_ VGND VGND VPWR VPWR _1247_ sky130_fd_sc_hd__or3_4
XFILLER_0_8_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4726_ _0707_ _3719_ _0100_ _0477_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4657_ _0024_ _0025_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__xor2_1
XFILLER_0_114_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7445_ _1045_ _1034_ _0925_ VGND VGND VPWR VPWR _3071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7376_ _1045_ net54 VGND VGND VPWR VPWR _2997_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4588_ _3688_ _3690_ VGND VGND VPWR VPWR _3691_ sky130_fd_sc_hd__or2_1
X_6327_ _1815_ _1849_ VGND VGND VPWR VPWR _1850_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6258_ _0829_ _1774_ _1000_ VGND VGND VPWR VPWR _1775_ sky130_fd_sc_hd__a21o_1
X_5209_ _0624_ _0627_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__xnor2_2
X_6189_ _1696_ _1697_ _1534_ _1536_ VGND VGND VPWR VPWR _1699_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3890_ net17 VGND VGND VPWR VPWR _1745_ sky130_fd_sc_hd__buf_2
XFILLER_0_57_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5560_ _1009_ _1010_ VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__or2_2
XFILLER_0_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4511_ _3521_ _3528_ VGND VGND VPWR VPWR _3614_ sky130_fd_sc_hd__or2b_1
XFILLER_0_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5491_ _3644_ _3619_ _0933_ _0934_ VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_14_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4442_ _3543_ _3544_ _3535_ VGND VGND VPWR VPWR _3546_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7230_ _2822_ _2823_ _2836_ _2837_ VGND VGND VPWR VPWR _2838_ sky130_fd_sc_hd__a211o_1
XFILLER_0_111_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4373_ _3476_ _3477_ _3384_ VGND VGND VPWR VPWR _3478_ sky130_fd_sc_hd__o21ai_1
X_7161_ _2739_ _2741_ _2760_ _2761_ VGND VGND VPWR VPWR _2763_ sky130_fd_sc_hd__nand4_4
XFILLER_0_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6112_ _1611_ _1614_ VGND VGND VPWR VPWR _1615_ sky130_fd_sc_hd__nand2_1
X_7092_ _1939_ _2687_ _0866_ VGND VGND VPWR VPWR _2688_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6043_ _1536_ _1538_ _1522_ VGND VGND VPWR VPWR _1540_ sky130_fd_sc_hd__a21oi_2
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6945_ _3273_ _1931_ _1952_ _3198_ VGND VGND VPWR VPWR _2526_ sky130_fd_sc_hd__a22oi_1
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6876_ _2450_ VGND VGND VPWR VPWR _2451_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5827_ _1299_ _1301_ VGND VGND VPWR VPWR _1303_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5758_ _0373_ net9 net10 _3352_ VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4709_ _3609_ _3682_ _0082_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7428_ _1603_ _1668_ _3052_ VGND VGND VPWR VPWR _3053_ sky130_fd_sc_hd__and3b_1
X_5689_ _1015_ _1016_ _1032_ _1152_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__a211o_2
XFILLER_0_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7359_ _3386_ _1963_ VGND VGND VPWR VPWR _2978_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4991_ _0253_ _0262_ _0261_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_81_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6730_ _3712_ _2278_ _2279_ _0309_ VGND VGND VPWR VPWR _2291_ sky130_fd_sc_hd__o22a_1
XFILLER_0_129_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3942_ _2302_ VGND VGND VPWR VPWR _2313_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3873_ _1373_ _1406_ _1537_ VGND VGND VPWR VPWR _1559_ sky130_fd_sc_hd__nand3_1
X_6661_ _2071_ _2080_ VGND VGND VPWR VPWR _2216_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6592_ _2136_ _2137_ _2139_ VGND VGND VPWR VPWR _2140_ sky130_fd_sc_hd__nand3_1
X_5612_ _0932_ _0940_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5543_ _0990_ _0992_ _0810_ _0896_ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__a211o_1
XFILLER_0_6_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5474_ _0905_ _0917_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_112_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4425_ _3521_ _3528_ VGND VGND VPWR VPWR _3529_ sky130_fd_sc_hd__xnor2_1
X_7213_ _2622_ _2818_ VGND VGND VPWR VPWR _2820_ sky130_fd_sc_hd__or2_1
X_4356_ _3356_ _3364_ _3363_ VGND VGND VPWR VPWR _3461_ sky130_fd_sc_hd__a21bo_1
X_7144_ _0174_ _2543_ _2576_ _3720_ VGND VGND VPWR VPWR _2744_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_1_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4287_ _3389_ _3391_ VGND VGND VPWR VPWR _3393_ sky130_fd_sc_hd__nand2_1
X_7075_ _2667_ _2668_ VGND VGND VPWR VPWR _2669_ sky130_fd_sc_hd__nor2_1
X_6026_ _1369_ _1377_ VGND VGND VPWR VPWR _1521_ sky130_fd_sc_hd__or2b_1
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6928_ _2504_ _2505_ _2506_ VGND VGND VPWR VPWR _2507_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6859_ _2419_ _2420_ _2430_ VGND VGND VPWR VPWR _2432_ sky130_fd_sc_hd__nand3_1
XFILLER_0_147_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4210_ _3242_ _3176_ net29 net30 VGND VGND VPWR VPWR _3317_ sky130_fd_sc_hd__nand4_2
XFILLER_0_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5190_ _0599_ _0606_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__xnor2_2
X_4141_ _3245_ _3246_ _3247_ VGND VGND VPWR VPWR _3249_ sky130_fd_sc_hd__a21o_1
X_4072_ _0270_ _1471_ _1460_ VGND VGND VPWR VPWR _3181_ sky130_fd_sc_hd__a21o_1
XFILLER_0_116_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4974_ _0042_ _2215_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3925_ _2117_ VGND VGND VPWR VPWR _2127_ sky130_fd_sc_hd__clkbuf_4
X_6713_ _2131_ _2272_ VGND VGND VPWR VPWR _2273_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_129_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6644_ _2027_ _2028_ _2047_ _2048_ VGND VGND VPWR VPWR _2197_ sky130_fd_sc_hd__a211o_2
XFILLER_0_144_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3856_ _1329_ _1362_ VGND VGND VPWR VPWR _1373_ sky130_fd_sc_hd__or2b_1
XFILLER_0_73_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3787_ _0150_ _0608_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6575_ _0855_ _1950_ _1951_ _0854_ _2121_ VGND VGND VPWR VPWR _2122_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5526_ _0972_ _0973_ _0974_ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__nand3_4
XFILLER_0_14_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5457_ _0723_ _0736_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4408_ _3511_ VGND VGND VPWR VPWR _3512_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5388_ _0820_ _0822_ _0819_ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4339_ _0030_ _2302_ _2368_ _3169_ VGND VGND VPWR VPWR _3444_ sky130_fd_sc_hd__a22o_1
X_7127_ _2722_ _2723_ _2724_ VGND VGND VPWR VPWR _2725_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7058_ _2647_ _2648_ _2612_ _2613_ VGND VGND VPWR VPWR _2650_ sky130_fd_sc_hd__o211ai_2
X_6009_ _3530_ _2117_ _0326_ _0453_ VGND VGND VPWR VPWR _1502_ sky130_fd_sc_hd__nand4_2
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_722 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4690_ _0040_ _0060_ _0061_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6360_ _1729_ _1724_ VGND VGND VPWR VPWR _1886_ sky130_fd_sc_hd__and2b_1
X_5311_ _0609_ _0611_ _0737_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__or3_1
XFILLER_0_12_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6291_ _1808_ _1809_ VGND VGND VPWR VPWR _1811_ sky130_fd_sc_hd__xnor2_2
X_5242_ _0664_ _0458_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__nor2_1
X_5173_ _0572_ _0578_ _0582_ _0589_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__a211o_1
X_4124_ net1 net60 _3172_ VGND VGND VPWR VPWR _3232_ sky130_fd_sc_hd__and3_1
Xinput1 A[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_4
X_4055_ _2914_ _3160_ _3162_ _3163_ VGND VGND VPWR VPWR _3164_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_94_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4957_ _0344_ _0352_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4888_ _0275_ _0276_ _0210_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__a21oi_1
X_3908_ _1931_ VGND VGND VPWR VPWR _1942_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3839_ _1165_ _1144_ _1154_ net65 VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__and4bb_2
X_6627_ _2176_ _2177_ VGND VGND VPWR VPWR _2178_ sky130_fd_sc_hd__or2b_1
XFILLER_0_34_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6558_ _2100_ _2101_ _1965_ net174 VGND VGND VPWR VPWR _2103_ sky130_fd_sc_hd__a211o_1
XFILLER_0_132_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5509_ _0948_ _0955_ VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__xor2_1
X_6489_ _1899_ _1900_ VGND VGND VPWR VPWR _2027_ sky130_fd_sc_hd__or2b_1
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_788 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5860_ _1174_ _1182_ VGND VGND VPWR VPWR _1339_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4811_ _0980_ _0870_ _0969_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__or3_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5791_ _1262_ _1263_ VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_75_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4742_ _0094_ _0096_ _0116_ _0118_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4673_ _0041_ _2106_ _2149_ _3645_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__a22oi_2
X_7461_ _0237_ _3158_ _1220_ VGND VGND VPWR VPWR _3088_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6412_ _0855_ _1928_ _1929_ _0854_ VGND VGND VPWR VPWR _1944_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7392_ _3012_ _3014_ VGND VGND VPWR VPWR _3015_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6343_ _1859_ _1860_ _1866_ VGND VGND VPWR VPWR _1868_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6274_ _1643_ _1644_ _1676_ _1677_ VGND VGND VPWR VPWR _1792_ sky130_fd_sc_hd__o211ai_2
X_5225_ _0519_ _0613_ _0644_ _0645_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_44_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5156_ net25 VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__buf_2
XFILLER_0_47_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4107_ _3202_ _3214_ VGND VGND VPWR VPWR _3215_ sky130_fd_sc_hd__nand2_2
X_5087_ _3388_ _0493_ _0494_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__and3_1
X_4038_ _1821_ _2007_ _2029_ VGND VGND VPWR VPWR _3147_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_614 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5989_ _1478_ _1479_ VGND VGND VPWR VPWR _1480_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_758 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5010_ _0279_ _0280_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__nand2_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6961_ _0100_ _2499_ _2543_ _3719_ VGND VGND VPWR VPWR _2544_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5912_ _3531_ net10 net11 _0161_ VGND VGND VPWR VPWR _1397_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6892_ _2453_ _2454_ _2466_ _2468_ VGND VGND VPWR VPWR _2469_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_146_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5843_ _1166_ _1167_ VGND VGND VPWR VPWR _1321_ sky130_fd_sc_hd__and2b_1
XFILLER_0_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5774_ _1241_ _1243_ _1244_ VGND VGND VPWR VPWR _1246_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_8_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4725_ _0099_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4656_ _3616_ _3618_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__or2_1
X_7444_ _0863_ _1067_ _3211_ VGND VGND VPWR VPWR _3070_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4587_ _3575_ _3577_ _3689_ VGND VGND VPWR VPWR _3690_ sky130_fd_sc_hd__a21o_1
X_7375_ _3209_ net57 VGND VGND VPWR VPWR _2996_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6326_ _1846_ _1847_ VGND VGND VPWR VPWR _1849_ sky130_fd_sc_hd__or2b_1
XFILLER_0_149_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6257_ _0693_ _0694_ _0830_ VGND VGND VPWR VPWR _1774_ sky130_fd_sc_hd__a21o_1
X_5208_ _0625_ _0626_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__nor2_1
X_6188_ _1534_ _1536_ _1696_ _1697_ VGND VGND VPWR VPWR _1698_ sky130_fd_sc_hd__a211oi_4
X_5139_ _0550_ _0551_ _0083_ _0170_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_99_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4510_ _3519_ _3552_ _3553_ VGND VGND VPWR VPWR _3613_ sky130_fd_sc_hd__nand3_2
X_5490_ _0933_ _0934_ _3644_ _3619_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_5_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4441_ _3535_ _3543_ _3544_ VGND VGND VPWR VPWR _3545_ sky130_fd_sc_hd__nand3_2
XFILLER_0_102_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7160_ _2758_ _2759_ _2553_ _2556_ VGND VGND VPWR VPWR _2761_ sky130_fd_sc_hd__o211ai_4
X_4372_ _3381_ _3475_ VGND VGND VPWR VPWR _3477_ sky130_fd_sc_hd__and2_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6111_ _1456_ _1305_ _1452_ _1612_ VGND VGND VPWR VPWR _1614_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7091_ _2018_ _2007_ _1821_ _1810_ _0863_ _0864_ VGND VGND VPWR VPWR _2687_ sky130_fd_sc_hd__mux4_1
X_6042_ _1522_ _1536_ _1538_ VGND VGND VPWR VPWR _1539_ sky130_fd_sc_hd__and3_2
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6944_ _2903_ _1952_ _2347_ _2345_ VGND VGND VPWR VPWR _2525_ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6875_ _2254_ _2243_ VGND VGND VPWR VPWR _2450_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5826_ _1299_ _1301_ VGND VGND VPWR VPWR _1302_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5757_ _3352_ _0373_ net9 VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4708_ _3610_ _3681_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5688_ _0320_ _1150_ _1151_ VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__and3_1
X_7427_ _0925_ _1067_ _3209_ _0969_ VGND VGND VPWR VPWR _3052_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4639_ _3414_ _3721_ _3722_ _3194_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7358_ _0063_ _1821_ VGND VGND VPWR VPWR _2977_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7289_ _1067_ net56 VGND VGND VPWR VPWR _2901_ sky130_fd_sc_hd__nand2_1
X_6309_ _1662_ _1664_ VGND VGND VPWR VPWR _1830_ sky130_fd_sc_hd__nand2_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4990_ _0386_ _0387_ _0377_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3941_ net28 VGND VGND VPWR VPWR _2302_ sky130_fd_sc_hd__buf_4
XFILLER_0_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3872_ _1373_ _1406_ _1537_ VGND VGND VPWR VPWR _1548_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6660_ _2079_ _2074_ VGND VGND VPWR VPWR _2214_ sky130_fd_sc_hd__or2b_1
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6591_ _1993_ _1994_ _1992_ VGND VGND VPWR VPWR _2139_ sky130_fd_sc_hd__a21bo_1
X_5611_ _0944_ _0945_ _0979_ _0981_ VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__nor4_1
XFILLER_0_6_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5542_ _0810_ _0896_ _0990_ _0992_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5473_ _0915_ _0916_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4424_ _3522_ _3527_ VGND VGND VPWR VPWR _3528_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7212_ _2622_ _2818_ VGND VGND VPWR VPWR _2819_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4355_ _3457_ _3458_ _3446_ VGND VGND VPWR VPWR _3460_ sky130_fd_sc_hd__a21o_1
X_7143_ _2524_ _2531_ VGND VGND VPWR VPWR _2743_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7074_ _2500_ _2497_ _2666_ _3192_ VGND VGND VPWR VPWR _2668_ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4286_ _3389_ _3391_ VGND VGND VPWR VPWR _3392_ sky130_fd_sc_hd__or2_1
X_6025_ _1375_ _1376_ VGND VGND VPWR VPWR _1520_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6927_ _0303_ net20 VGND VGND VPWR VPWR _2506_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6858_ _2419_ _2420_ _2430_ VGND VGND VPWR VPWR _2431_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5809_ _0710_ _1283_ _0429_ VGND VGND VPWR VPWR _1284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6789_ _2155_ _2157_ VGND VGND VPWR VPWR _2355_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4140_ _3245_ _3246_ _3247_ VGND VGND VPWR VPWR _3248_ sky130_fd_sc_hd__nand3_1
X_4071_ _3177_ _3178_ _3175_ VGND VGND VPWR VPWR _3180_ sky130_fd_sc_hd__a21o_1
XFILLER_0_116_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4973_ _0369_ _0370_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3924_ _2106_ VGND VGND VPWR VPWR _2117_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6712_ _2268_ _2271_ VGND VGND VPWR VPWR _2272_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6643_ net143 VGND VGND VPWR VPWR _2196_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3855_ _0980_ _1002_ _1340_ _1351_ VGND VGND VPWR VPWR _1362_ sky130_fd_sc_hd__a31o_1
XFILLER_0_74_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3786_ _0259_ _0576_ _0597_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__a21o_1
X_6574_ _0199_ _0428_ _3707_ _3161_ VGND VGND VPWR VPWR _2121_ sky130_fd_sc_hd__o31a_1
XFILLER_0_144_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5525_ _0784_ _0792_ _0791_ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_14_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5456_ _0734_ _0735_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4407_ net34 VGND VGND VPWR VPWR _3511_ sky130_fd_sc_hd__clkbuf_4
X_5387_ _0819_ _0820_ _0822_ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4338_ _3169_ net191 _2302_ VGND VGND VPWR VPWR _3443_ sky130_fd_sc_hd__and3_1
X_7126_ _2512_ _2517_ _2511_ VGND VGND VPWR VPWR _2724_ sky130_fd_sc_hd__a21bo_1
X_4269_ _3372_ _3373_ _3340_ VGND VGND VPWR VPWR _3375_ sky130_fd_sc_hd__o21ai_2
X_7057_ _2612_ _2613_ _2647_ _2648_ VGND VGND VPWR VPWR _2649_ sky130_fd_sc_hd__a211o_1
X_6008_ _2117_ _0219_ _1366_ _1365_ VGND VGND VPWR VPWR _1501_ sky130_fd_sc_hd__a31o_1
XFILLER_0_69_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5310_ _0609_ _0611_ _0737_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_12_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6290_ _1631_ _1634_ VGND VGND VPWR VPWR _1809_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5241_ _0445_ _0991_ _0327_ _0454_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__and4_1
X_5172_ _0428_ _0586_ _0588_ _0849_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4123_ _1439_ _3186_ _3187_ VGND VGND VPWR VPWR _3231_ sky130_fd_sc_hd__nand3b_1
Xinput2 A[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_4
X_4054_ _0925_ _0969_ _1100_ VGND VGND VPWR VPWR _3163_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4956_ _0350_ _0351_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4887_ _0210_ _0275_ _0276_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__and3_1
XFILLER_0_117_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3907_ net15 VGND VGND VPWR VPWR _1931_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_117_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3838_ _0783_ _1144_ _1154_ _1165_ VGND VGND VPWR VPWR _1176_ sky130_fd_sc_hd__nor4b_2
X_6626_ _3512_ _2532_ _2565_ _3423_ VGND VGND VPWR VPWR _2177_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6557_ _1965_ net175 _2100_ net171 VGND VGND VPWR VPWR _2102_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_132_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5508_ _0949_ _0954_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__xnor2_1
X_3769_ _0412_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__buf_2
XFILLER_0_15_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6488_ _2023_ _2024_ _1870_ _1991_ VGND VGND VPWR VPWR _2026_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5439_ _0826_ _0836_ _0878_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__o21bai_1
X_7109_ _2353_ _2503_ _2534_ _2535_ VGND VGND VPWR VPWR _2705_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4810_ net124 _0175_ _3204_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5790_ _1132_ _1135_ VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__or2b_4
XFILLER_0_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4741_ _0097_ _0098_ _0115_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4672_ _0042_ _3530_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__nand2_1
X_7460_ _1613_ _1635_ _1668_ VGND VGND VPWR VPWR _3086_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6411_ _0848_ _1940_ _1941_ _0849_ VGND VGND VPWR VPWR _1943_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7391_ _3486_ _2007_ VGND VGND VPWR VPWR _3014_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6342_ _1859_ _1860_ _1866_ VGND VGND VPWR VPWR _1867_ sky130_fd_sc_hd__nand3_1
XFILLER_0_12_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6273_ _1475_ _1637_ VGND VGND VPWR VPWR _1791_ sky130_fd_sc_hd__nand2_1
X_5224_ _0642_ _0643_ _0623_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__a21oi_2
X_5155_ _0439_ _0425_ _0563_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4106_ _2401_ _3198_ VGND VGND VPWR VPWR _3214_ sky130_fd_sc_hd__nand2_1
X_5086_ _3433_ _3431_ net32 net2 VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__nand4_2
XFILLER_0_47_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4037_ _1767_ _1799_ _0892_ VGND VGND VPWR VPWR _3146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5988_ _1355_ _1357_ _1477_ VGND VGND VPWR VPWR _1479_ sky130_fd_sc_hd__or3_1
X_4939_ _0222_ _0230_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__or2b_1
XFILLER_0_93_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_636 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6609_ _3385_ _2609_ _2155_ _2156_ VGND VGND VPWR VPWR _2158_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_34_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_718 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_306 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_578 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6960_ _3719_ _0100_ _2499_ VGND VGND VPWR VPWR _2542_ sky130_fd_sc_hd__and3_1
X_5911_ _0161_ _0373_ _2565_ VGND VGND VPWR VPWR _1396_ sky130_fd_sc_hd__and3_1
X_6891_ _2455_ _2211_ _2465_ VGND VGND VPWR VPWR _2468_ sky130_fd_sc_hd__and3_1
XFILLER_0_124_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5842_ _1189_ _1191_ VGND VGND VPWR VPWR _1320_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5773_ _1241_ _1243_ _1244_ VGND VGND VPWR VPWR _1245_ sky130_fd_sc_hd__and3_2
XFILLER_0_75_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4724_ net37 VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4655_ _0022_ _0023_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__nor2_1
X_7443_ _3065_ _3067_ _3068_ VGND VGND VPWR VPWR _3069_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7374_ _2739_ _2763_ VGND VGND VPWR VPWR _2995_ sky130_fd_sc_hd__nand2_1
X_4586_ _3513_ _2237_ VGND VGND VPWR VPWR _3689_ sky130_fd_sc_hd__and2b_1
Xinput60 B[5] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6325_ _1815_ _1846_ _1847_ VGND VGND VPWR VPWR _1848_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_101_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6256_ _1448_ VGND VGND VPWR VPWR _1773_ sky130_fd_sc_hd__inv_2
X_5207_ _3645_ _0041_ _2686_ _2740_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__and4_1
X_6187_ _1694_ _1695_ _1681_ VGND VGND VPWR VPWR _1697_ sky130_fd_sc_hd__a21oi_2
X_5138_ _0286_ _0415_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5069_ _3442_ _2434_ _0104_ _3511_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__nand4_2
XFILLER_0_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4440_ _3540_ _3541_ _3542_ VGND VGND VPWR VPWR _3544_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4371_ _3381_ _3475_ VGND VGND VPWR VPWR _3476_ sky130_fd_sc_hd__nor2_2
XFILLER_0_0_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6110_ _1297_ _1450_ _1451_ VGND VGND VPWR VPWR _1612_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_95_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7090_ _0854_ _2670_ _2671_ _0855_ _2684_ VGND VGND VPWR VPWR _2685_ sky130_fd_sc_hd__a221o_1
X_6041_ _1534_ _1535_ _1528_ VGND VGND VPWR VPWR _1538_ sky130_fd_sc_hd__a21o_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6943_ _2358_ _2360_ VGND VGND VPWR VPWR _2524_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6874_ _1067_ _1384_ _2263_ _2299_ VGND VGND VPWR VPWR _2449_ sky130_fd_sc_hd__and4_2
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5825_ _1272_ _1274_ _1300_ VGND VGND VPWR VPWR _1301_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5756_ _1217_ _1225_ VGND VGND VPWR VPWR _1226_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4707_ _0079_ _0080_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__nor2_1
X_5687_ _1146_ _1149_ _1142_ VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7426_ _0860_ _0712_ VGND VGND VPWR VPWR _3051_ sky130_fd_sc_hd__nor2_1
X_4638_ _3580_ _3118_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4569_ _3517_ _3670_ _3671_ VGND VGND VPWR VPWR _3672_ sky130_fd_sc_hd__nor3_4
X_7357_ _2710_ _2712_ VGND VGND VPWR VPWR _2976_ sky130_fd_sc_hd__nand2_1
X_7288_ _2863_ _2865_ _2860_ VGND VGND VPWR VPWR _2900_ sky130_fd_sc_hd__o21ai_1
X_6308_ _1820_ _1828_ VGND VGND VPWR VPWR _1829_ sky130_fd_sc_hd__xor2_1
X_6239_ _1626_ _1753_ VGND VGND VPWR VPWR _1754_ sky130_fd_sc_hd__xor2_2
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_670 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3940_ _2193_ _2281_ _0936_ VGND VGND VPWR VPWR _2292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3871_ _1515_ _1526_ VGND VGND VPWR VPWR _1537_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6590_ _2133_ _2134_ _2135_ VGND VGND VPWR VPWR _2137_ sky130_fd_sc_hd__a21o_1
X_5610_ _1063_ _1064_ _1037_ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5541_ _0988_ _0989_ _0897_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5472_ _0724_ _0732_ _0731_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__a21bo_1
X_7211_ _2815_ _2816_ VGND VGND VPWR VPWR _2818_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4423_ _3525_ _3526_ VGND VGND VPWR VPWR _3527_ sky130_fd_sc_hd__or2_2
XFILLER_0_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4354_ _3446_ _3457_ _3458_ VGND VGND VPWR VPWR _3459_ sky130_fd_sc_hd__nand3_2
X_7142_ _2525_ _2530_ VGND VGND VPWR VPWR _2742_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7073_ _2500_ _2497_ _2666_ VGND VGND VPWR VPWR _2667_ sky130_fd_sc_hd__a21oi_1
X_4285_ _3276_ _3278_ _3390_ VGND VGND VPWR VPWR _3391_ sky130_fd_sc_hd__a21o_1
X_6024_ _1516_ _1517_ _1350_ _1481_ VGND VGND VPWR VPWR _1519_ sky130_fd_sc_hd__a211o_1
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6926_ _0881_ _0521_ net21 net22 VGND VGND VPWR VPWR _2505_ sky130_fd_sc_hd__nand4_2
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6857_ _2421_ _2429_ VGND VGND VPWR VPWR _2430_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6788_ _2350_ _2351_ _2352_ VGND VGND VPWR VPWR _2354_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5808_ _1909_ _1876_ _0862_ _2587_ _0583_ _0584_ VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__mux4_1
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5739_ _1205_ _1206_ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_745 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7409_ _3031_ _3032_ VGND VGND VPWR VPWR _3033_ sky130_fd_sc_hd__xnor2_1
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4070_ _3175_ _3177_ net195 VGND VGND VPWR VPWR _3179_ sky130_fd_sc_hd__nand3_1
XFILLER_0_116_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4972_ _0366_ _0367_ _0360_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3923_ net31 VGND VGND VPWR VPWR _2106_ sky130_fd_sc_hd__buf_4
XFILLER_0_86_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6711_ _2269_ net170 VGND VGND VPWR VPWR _2271_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3854_ _0881_ _0357_ _0717_ VGND VGND VPWR VPWR _1351_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6642_ _2070_ _2082_ _2083_ VGND VGND VPWR VPWR _2195_ sky130_fd_sc_hd__and3_1
XFILLER_0_144_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3785_ _0587_ _0226_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6573_ _0438_ _2119_ _1277_ VGND VGND VPWR VPWR _2120_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5524_ _0970_ _0971_ _0962_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5455_ _0738_ _0742_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4406_ _3428_ _3438_ VGND VGND VPWR VPWR _3510_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5386_ _0549_ _0552_ _0553_ _0821_ VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__a31o_1
X_7125_ _2714_ _2715_ _2721_ VGND VGND VPWR VPWR _2723_ sky130_fd_sc_hd__a21o_1
X_4337_ net29 VGND VGND VPWR VPWR _3442_ sky130_fd_sc_hd__buf_4
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4268_ _3340_ _3372_ _3373_ VGND VGND VPWR VPWR _3374_ sky130_fd_sc_hd__or3_4
X_7056_ _2645_ _2646_ _2436_ _2438_ VGND VGND VPWR VPWR _2648_ sky130_fd_sc_hd__o211a_1
X_6007_ _1342_ _1344_ VGND VGND VPWR VPWR _1500_ sky130_fd_sc_hd__or2_1
X_4199_ _3236_ _3239_ _3237_ VGND VGND VPWR VPWR _3306_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_96_326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6909_ _2327_ _2328_ _2485_ _2486_ VGND VGND VPWR VPWR _2487_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_147_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_779 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5240_ _0660_ _0661_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5171_ _3210_ _0196_ _3727_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4122_ _3218_ _3229_ VGND VGND VPWR VPWR _3230_ sky130_fd_sc_hd__or2b_1
X_4053_ _0870_ _0063_ _3161_ VGND VGND VPWR VPWR _3162_ sky130_fd_sc_hd__and3_2
Xinput3 A[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_4
XFILLER_0_127_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4955_ _0224_ _0225_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3906_ _1876_ _1909_ _0892_ VGND VGND VPWR VPWR _1920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4886_ _0273_ _0274_ _0153_ _0155_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__a211o_1
XFILLER_0_7_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3837_ net66 VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__clkbuf_2
X_6625_ _3423_ _3512_ _2532_ _2565_ VGND VGND VPWR VPWR _2176_ sky130_fd_sc_hd__and4_1
XFILLER_0_7_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3768_ net12 VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__buf_6
XFILLER_0_61_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6556_ _2098_ _2099_ _1966_ _1967_ VGND VGND VPWR VPWR _2101_ sky130_fd_sc_hd__a211o_1
XFILLER_0_131_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5507_ _0952_ _0953_ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6487_ _1870_ _1991_ _2023_ _2024_ VGND VGND VPWR VPWR _2025_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5438_ _0876_ _0877_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__or2_2
XFILLER_0_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5369_ _0766_ _0767_ _0801_ _0802_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__nor4_4
XFILLER_0_100_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7108_ _2564_ _2566_ _2605_ _2606_ VGND VGND VPWR VPWR _2704_ sky130_fd_sc_hd__and4bb_1
X_7039_ _2402_ _2405_ VGND VGND VPWR VPWR _2629_ sky130_fd_sc_hd__or2_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_749 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4740_ _0097_ _0098_ _0115_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4671_ net60 VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7390_ _3007_ _3011_ VGND VGND VPWR VPWR _3012_ sky130_fd_sc_hd__xnor2_1
X_6410_ _0848_ _3503_ VGND VGND VPWR VPWR _1941_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6341_ _1863_ _1864_ VGND VGND VPWR VPWR _1866_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6272_ _1743_ VGND VGND VPWR VPWR _1790_ sky130_fd_sc_hd__inv_2
X_5223_ _0623_ _0642_ _0643_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5154_ _0439_ _0425_ _0563_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__nand3_1
XFILLER_0_138_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4105_ _3207_ _3212_ _1100_ VGND VGND VPWR VPWR _3213_ sky130_fd_sc_hd__mux2_2
X_5085_ net162 net32 net2 net61 VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__a22o_4
X_4036_ _3143_ _3144_ _3131_ VGND VGND VPWR VPWR _3145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5987_ _1355_ _1357_ _1477_ VGND VGND VPWR VPWR _1478_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4938_ _0225_ _0227_ _0229_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__or3_2
X_4869_ _0254_ _0255_ _0256_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__nand3_1
XFILLER_0_62_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6608_ _2155_ _2156_ _3385_ _2598_ VGND VGND VPWR VPWR _2157_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_7_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6539_ _1836_ _1838_ _2081_ VGND VGND VPWR VPWR _2082_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_638 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5910_ _1385_ _1393_ VGND VGND VPWR VPWR _1394_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6890_ _2455_ _2211_ _2465_ VGND VGND VPWR VPWR _2466_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_124_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5841_ _1317_ VGND VGND VPWR VPWR _1319_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5772_ _1106_ _1115_ _1114_ VGND VGND VPWR VPWR _1244_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_57_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4723_ _0032_ _0039_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7442_ _1165_ _0783_ _1144_ _1154_ VGND VGND VPWR VPWR _3068_ sky130_fd_sc_hd__or4b_1
XFILLER_0_140_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4654_ _0423_ _3619_ _0020_ _0021_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_71_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7373_ _2748_ _2756_ _2993_ VGND VGND VPWR VPWR _2994_ sky130_fd_sc_hd__o21ai_1
X_4585_ _3686_ _3687_ VGND VGND VPWR VPWR _3688_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput61 B[6] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_8
Xinput50 B[25] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_114_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6324_ _1844_ _1845_ _1696_ _1698_ VGND VGND VPWR VPWR _1847_ sky130_fd_sc_hd__a211o_1
XFILLER_0_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6255_ _0563_ _0693_ _0829_ _0878_ VGND VGND VPWR VPWR _1772_ sky130_fd_sc_hd__and4_1
X_5206_ _0041_ _2696_ _2740_ _0172_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__a22oi_2
X_6186_ _1681_ _1694_ _1695_ VGND VGND VPWR VPWR _1696_ sky130_fd_sc_hd__and3_2
X_5137_ _0081_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__inv_2
X_5068_ _2423_ _3422_ _3511_ _2368_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__a22o_1
X_4019_ _2543_ VGND VGND VPWR VPWR _3128_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_109_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4370_ _3472_ _3474_ VGND VGND VPWR VPWR _3475_ sky130_fd_sc_hd__xor2_1
XFILLER_0_111_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6040_ _1528_ _1534_ _1535_ VGND VGND VPWR VPWR _1536_ sky130_fd_sc_hd__nand3_2
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6942_ _2518_ _2519_ _2520_ VGND VGND VPWR VPWR _2523_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_49_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6873_ _1067_ _2263_ _2299_ _3209_ VGND VGND VPWR VPWR _2448_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_146_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5824_ _1170_ _1909_ VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__and2b_1
XFILLER_0_146_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5755_ _1218_ _1224_ VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4706_ _3679_ _0078_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__and2_1
X_5686_ _1142_ _1146_ _1149_ VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__nand3_1
XFILLER_0_97_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7425_ _3127_ _0703_ _3049_ VGND VGND VPWR VPWR _3050_ sky130_fd_sc_hd__a21o_1
X_4637_ _0003_ _0005_ _3301_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4568_ _3668_ _3669_ _3552_ _3613_ VGND VGND VPWR VPWR _3671_ sky130_fd_sc_hd__o211a_1
X_7356_ _2903_ _1778_ _2719_ _2717_ VGND VGND VPWR VPWR _2975_ sky130_fd_sc_hd__a31o_1
XFILLER_0_69_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4499_ _3207_ _3602_ _3077_ VGND VGND VPWR VPWR _3603_ sky130_fd_sc_hd__mux2_1
X_6307_ _1826_ _1827_ VGND VGND VPWR VPWR _1828_ sky130_fd_sc_hd__nand2_1
X_7287_ _3144_ _0196_ _2319_ _2894_ _2898_ VGND VGND VPWR VPWR _2899_ sky130_fd_sc_hd__o311a_1
X_6238_ _1628_ _1752_ VGND VGND VPWR VPWR _1753_ sky130_fd_sc_hd__xor2_4
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _1674_ _1675_ _1539_ _1541_ VGND VGND VPWR VPWR _1677_ sky130_fd_sc_hd__a211o_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3870_ _1417_ _1439_ _1504_ VGND VGND VPWR VPWR _1526_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5540_ _0897_ _0988_ _0989_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5471_ _0906_ _0913_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_724 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4422_ _0324_ _3343_ _3523_ _3524_ VGND VGND VPWR VPWR _3526_ sky130_fd_sc_hd__and4_1
XFILLER_0_30_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7210_ _3209_ net56 VGND VGND VPWR VPWR _2816_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4353_ _3454_ _3455_ _3456_ VGND VGND VPWR VPWR _3458_ sky130_fd_sc_hd__a21o_1
X_7141_ _2737_ _2738_ _2522_ _2708_ VGND VGND VPWR VPWR _2741_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4284_ _3273_ _3139_ VGND VGND VPWR VPWR _3390_ sky130_fd_sc_hd__and2b_1
X_7072_ _2663_ _2665_ VGND VGND VPWR VPWR _2666_ sky130_fd_sc_hd__or2_1
X_6023_ _1350_ _1481_ _1516_ _1517_ VGND VGND VPWR VPWR _1518_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_146_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6925_ _0521_ net21 net22 _0881_ VGND VGND VPWR VPWR _2504_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6856_ _2427_ _2428_ VGND VGND VPWR VPWR _2429_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3999_ _2914_ _2925_ VGND VGND VPWR VPWR _2936_ sky130_fd_sc_hd__or2_1
X_6787_ _2350_ _2351_ _2352_ VGND VGND VPWR VPWR _2353_ sky130_fd_sc_hd__and3_2
XFILLER_0_71_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5807_ _1270_ _1278_ _1279_ _1280_ _1281_ VGND VGND VPWR VPWR _1282_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_29_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5738_ _2215_ _0110_ VGND VGND VPWR VPWR _1206_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5669_ _1065_ _1066_ _1128_ _1129_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7408_ _2853_ _2855_ _2852_ VGND VGND VPWR VPWR _3032_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7339_ _2951_ _2955_ VGND VGND VPWR VPWR _2956_ sky130_fd_sc_hd__xnor2_1
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_608 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4971_ _0360_ _0366_ _0367_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3922_ _0870_ _1996_ _2084_ VGND VGND VPWR VPWR _2095_ sky130_fd_sc_hd__o21a_2
XFILLER_0_73_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6710_ _2093_ VGND VGND VPWR VPWR _2269_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3853_ _0881_ _0357_ _0717_ VGND VGND VPWR VPWR _1340_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6641_ _2082_ VGND VGND VPWR VPWR _2194_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3784_ _0172_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6572_ _1810_ _1949_ VGND VGND VPWR VPWR _2119_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5523_ _0962_ _0970_ _0971_ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__nand3_2
XFILLER_0_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5454_ _0719_ _0810_ _0811_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__nor3_1
XFILLER_0_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5385_ _0544_ _0545_ _0684_ VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__or3_4
X_4405_ _3437_ _3429_ VGND VGND VPWR VPWR _3509_ sky130_fd_sc_hd__and2b_1
X_4336_ _3440_ _2881_ VGND VGND VPWR VPWR _3441_ sky130_fd_sc_hd__nand2_1
X_7124_ _2714_ _2715_ _2721_ VGND VGND VPWR VPWR _2722_ sky130_fd_sc_hd__nand3_1
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4267_ _3370_ _3371_ _3327_ _3329_ VGND VGND VPWR VPWR _3373_ sky130_fd_sc_hd__o211a_1
X_7055_ _2436_ _2438_ _2645_ _2646_ VGND VGND VPWR VPWR _2647_ sky130_fd_sc_hd__a211oi_2
X_4198_ _1668_ VGND VGND VPWR VPWR _3305_ sky130_fd_sc_hd__buf_4
X_6006_ _1341_ _1348_ VGND VGND VPWR VPWR _1499_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_530 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6908_ _2483_ _2484_ _2329_ _2330_ VGND VGND VPWR VPWR _2486_ sky130_fd_sc_hd__a211o_1
XFILLER_0_108_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6839_ _2127_ _1007_ _2407_ _2408_ VGND VGND VPWR VPWR _2410_ sky130_fd_sc_hd__and4_1
XFILLER_0_147_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5170_ _1078_ _3407_ _0004_ _0585_ _0429_ _0189_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__mux4_1
X_4121_ _0063_ _3223_ _3228_ _3156_ VGND VGND VPWR VPWR _3229_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_127_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4052_ net25 net65 _1701_ VGND VGND VPWR VPWR _3161_ sky130_fd_sc_hd__and3_4
Xinput4 A[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4954_ _0345_ _0349_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__xor2_2
XFILLER_0_19_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3905_ _1898_ VGND VGND VPWR VPWR _1909_ sky130_fd_sc_hd__buf_4
XFILLER_0_74_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4885_ _0153_ net116 _0273_ _0274_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_62_717 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3836_ net68 VGND VGND VPWR VPWR _1154_ sky130_fd_sc_hd__clkbuf_2
X_6624_ _2173_ _2174_ VGND VGND VPWR VPWR _2175_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3767_ _0390_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__buf_4
XFILLER_0_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6555_ _1966_ _1967_ net157 _2099_ VGND VGND VPWR VPWR _2100_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_131_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5506_ _3343_ _2248_ _0950_ _0951_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__and4_1
XFILLER_0_14_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6486_ _2011_ _2012_ _2022_ VGND VGND VPWR VPWR _2024_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_30_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5437_ _0862_ _0875_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__and2_2
XFILLER_0_30_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5368_ _0799_ _0800_ _0642_ _0768_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4319_ _3423_ VGND VGND VPWR VPWR _3424_ sky130_fd_sc_hd__buf_4
X_5299_ _0194_ _0325_ _0452_ _0324_ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__a22oi_1
X_7107_ _2678_ _2701_ _2697_ VGND VGND VPWR VPWR _2703_ sky130_fd_sc_hd__a21o_1
X_7038_ _2459_ _2461_ VGND VGND VPWR VPWR _2628_ sky130_fd_sc_hd__or2_2
XFILLER_0_97_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_831 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4670_ _0032_ _0039_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__xor2_2
XFILLER_0_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6340_ _0042_ _1854_ VGND VGND VPWR VPWR _1864_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6271_ _1628_ _1752_ VGND VGND VPWR VPWR _1789_ sky130_fd_sc_hd__nand2_2
XFILLER_0_121_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5222_ _0638_ _0639_ _0640_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5153_ _0563_ _0567_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__xor2_1
X_4104_ _3208_ _3211_ _3131_ VGND VGND VPWR VPWR _3212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5084_ net60 _2204_ _0375_ _0374_ _0491_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__a32oi_2
X_4035_ _0903_ net25 VGND VGND VPWR VPWR _3144_ sky130_fd_sc_hd__or2b_2
XFILLER_0_79_647 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5986_ _1326_ _1327_ _1337_ _1475_ _1476_ VGND VGND VPWR VPWR _1477_ sky130_fd_sc_hd__o32ai_4
X_4937_ _0322_ _0330_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_20 net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4868_ _3449_ _3448_ _2686_ net6 VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__nand4_2
XFILLER_0_75_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6607_ _3272_ _1854_ _1898_ _3196_ VGND VGND VPWR VPWR _2156_ sky130_fd_sc_hd__a22oi_1
X_3819_ _0958_ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4799_ _3265_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_761 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6538_ _2071_ _2080_ VGND VGND VPWR VPWR _2081_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6469_ _2003_ _2004_ VGND VGND VPWR VPWR _2005_ sky130_fd_sc_hd__xor2_1
XFILLER_0_100_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5840_ _0904_ _1043_ _1156_ VGND VGND VPWR VPWR _1317_ sky130_fd_sc_hd__or3_1
XFILLER_0_124_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5771_ _1239_ _1240_ _1232_ VGND VGND VPWR VPWR _1243_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4722_ _0033_ _0038_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__or2b_1
XFILLER_0_57_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7441_ net57 _0571_ VGND VGND VPWR VPWR _3067_ sky130_fd_sc_hd__or2b_1
XFILLER_0_140_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4653_ _0020_ _0021_ _0423_ net35 VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__and4bb_1
Xinput40 B[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_2
XFILLER_0_142_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput51 B[26] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_4
X_7372_ _2754_ _2755_ VGND VGND VPWR VPWR _2993_ sky130_fd_sc_hd__nand2_1
X_4584_ _3137_ _3685_ VGND VGND VPWR VPWR _3687_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput62 B[7] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_6
XFILLER_0_40_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6323_ _1696_ _1698_ _1844_ _1845_ VGND VGND VPWR VPWR _1846_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6254_ _1011_ _1272_ _1299_ _1454_ VGND VGND VPWR VPWR _1771_ sky130_fd_sc_hd__and4_1
X_5205_ _0042_ _2653_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6185_ _1692_ _1693_ _1686_ VGND VGND VPWR VPWR _1695_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5136_ _0416_ _0547_ _0548_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_99_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5067_ _0471_ _0472_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__xnor2_2
X_4018_ _0063_ VGND VGND VPWR VPWR _3127_ sky130_fd_sc_hd__buf_2
XFILLER_0_95_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5969_ _1452_ _1457_ VGND VGND VPWR VPWR _1458_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6941_ _2518_ _2519_ _2520_ VGND VGND VPWR VPWR _2522_ sky130_fd_sc_hd__and3_2
XFILLER_0_44_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6872_ _3209_ _2263_ _2262_ VGND VGND VPWR VPWR _2447_ sky130_fd_sc_hd__nand3_1
XFILLER_0_44_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5823_ _1297_ _1298_ VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__or2_2
XFILLER_0_91_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5754_ _1222_ _1223_ VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4705_ _3679_ _0078_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__nor2_1
X_5685_ _0995_ _1147_ _1143_ _0820_ _1148_ VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__o221a_1
XFILLER_0_45_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7424_ _3162_ _3487_ _3048_ _0838_ VGND VGND VPWR VPWR _3049_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4636_ _3407_ _0004_ _3087_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7355_ _2970_ _2973_ VGND VGND VPWR VPWR _2974_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4567_ _3552_ _3613_ _3668_ _3669_ VGND VGND VPWR VPWR _3670_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_69_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6306_ _1824_ _1825_ _1651_ _1653_ VGND VGND VPWR VPWR _1827_ sky130_fd_sc_hd__a211o_1
X_4498_ _2237_ _2182_ _2138_ _3139_ _0925_ _0969_ VGND VGND VPWR VPWR _3602_ sky130_fd_sc_hd__mux4_1
XFILLER_0_13_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7286_ _2895_ _2896_ _2897_ VGND VGND VPWR VPWR _2898_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6237_ _1750_ _1751_ VGND VGND VPWR VPWR _1752_ sky130_fd_sc_hd__nor2_2
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _1539_ _1541_ _1674_ _1675_ VGND VGND VPWR VPWR _1676_ sky130_fd_sc_hd__o211ai_4
X_5119_ _0464_ _0528_ _0529_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__nand3_2
XFILLER_0_85_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6099_ _1138_ _1265_ _1434_ VGND VGND VPWR VPWR _1601_ sky130_fd_sc_hd__or3_1
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_560 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_472 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5470_ _0911_ _0912_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4421_ _0739_ _3430_ _3523_ _3524_ VGND VGND VPWR VPWR _3525_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_53_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4352_ _3454_ _3455_ _3456_ VGND VGND VPWR VPWR _3457_ sky130_fd_sc_hd__nand3_1
XFILLER_0_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7140_ _2522_ _2708_ _2737_ _2738_ VGND VGND VPWR VPWR _2739_ sky130_fd_sc_hd__o211ai_4
X_4283_ _3387_ _3388_ VGND VGND VPWR VPWR _3389_ sky130_fd_sc_hd__or2_2
X_7071_ _2501_ _2662_ VGND VGND VPWR VPWR _2665_ sky130_fd_sc_hd__and2_1
X_6022_ _1513_ _1514_ _1379_ _1381_ VGND VGND VPWR VPWR _1517_ sky130_fd_sc_hd__a211o_1
XFILLER_0_146_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6924_ _2353_ _2354_ _2365_ VGND VGND VPWR VPWR _2503_ sky130_fd_sc_hd__nor3_1
XFILLER_0_76_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6855_ _2425_ _2426_ _2172_ _2174_ VGND VGND VPWR VPWR _2428_ sky130_fd_sc_hd__o211ai_1
X_3998_ _2302_ net60 VGND VGND VPWR VPWR _2925_ sky130_fd_sc_hd__and2_2
XFILLER_0_91_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6786_ _2141_ _2146_ _2140_ VGND VGND VPWR VPWR _2352_ sky130_fd_sc_hd__a21bo_1
X_5806_ _0848_ _3097_ _3126_ VGND VGND VPWR VPWR _1281_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5737_ _1203_ _1204_ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__or2b_1
XFILLER_0_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5668_ _1065_ _1066_ _1128_ _1129_ VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__or4_4
XFILLER_0_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7407_ _2815_ _2816_ _2813_ VGND VGND VPWR VPWR _3031_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_32_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4619_ _2675_ _3720_ VGND VGND VPWR VPWR _3721_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5599_ _0929_ _0930_ _1052_ _1053_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__a211o_1
XFILLER_0_13_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7338_ _2952_ _2954_ VGND VGND VPWR VPWR _2955_ sky130_fd_sc_hd__xnor2_1
X_7269_ _0419_ _2699_ _2700_ _2879_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__a31o_4
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4970_ _0364_ _0365_ _0361_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3921_ _0554_ _2073_ _0587_ VGND VGND VPWR VPWR _2084_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3852_ _1307_ _1318_ VGND VGND VPWR VPWR _1329_ sky130_fd_sc_hd__xnor2_1
X_6640_ _2189_ _2190_ net189 net104 VGND VGND VPWR VPWR _2192_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_58_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_642 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6571_ _0861_ _2115_ _2116_ _0844_ VGND VGND VPWR VPWR _2118_ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5522_ _0966_ _0967_ _0968_ VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__a21o_1
X_3783_ _0379_ _0543_ _0565_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5453_ net140 net208 _0817_ _0682_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__and4b_1
X_5384_ _0540_ _0681_ _0684_ _0592_ VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__o22a_1
X_4404_ _1384_ _3425_ _3421_ VGND VGND VPWR VPWR _3508_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4335_ net194 VGND VGND VPWR VPWR _3440_ sky130_fd_sc_hd__clkbuf_4
X_7123_ _2719_ _2720_ VGND VGND VPWR VPWR _2721_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4266_ _3327_ _3329_ _3370_ net184 VGND VGND VPWR VPWR _3372_ sky130_fd_sc_hd__a211oi_2
X_7054_ _2643_ _2644_ _2624_ VGND VGND VPWR VPWR _2646_ sky130_fd_sc_hd__o21a_1
X_4197_ _2980_ _3282_ _3289_ _3303_ VGND VGND VPWR VPWR _3304_ sky130_fd_sc_hd__a211o_1
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6005_ _1488_ _1497_ VGND VGND VPWR VPWR _1498_ sky130_fd_sc_hd__xor2_2
XFILLER_0_77_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6907_ _2329_ _2330_ _2483_ _2484_ VGND VGND VPWR VPWR _2485_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_147_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6838_ _2127_ _1008_ _2407_ _2408_ VGND VGND VPWR VPWR _2409_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_147_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6769_ _2011_ _2132_ _2163_ _2164_ VGND VGND VPWR VPWR _2333_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_116_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4120_ _3200_ _3154_ _3227_ VGND VGND VPWR VPWR _3228_ sky130_fd_sc_hd__or3b_2
XFILLER_0_127_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4051_ _3158_ _3159_ _1220_ VGND VGND VPWR VPWR _3160_ sky130_fd_sc_hd__a21oi_1
Xinput5 A[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_4
XFILLER_0_36_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4953_ _3423_ _0347_ _0348_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_52_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3904_ _1887_ VGND VGND VPWR VPWR _1898_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4884_ _0234_ _0235_ _0271_ _0272_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_74_556 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6623_ _2718_ _0293_ _2170_ _2172_ VGND VGND VPWR VPWR _2174_ sky130_fd_sc_hd__nand4_2
XFILLER_0_52_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3835_ net67 VGND VGND VPWR VPWR _1144_ sky130_fd_sc_hd__buf_2
XFILLER_0_74_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3766_ net44 VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6554_ net169 _2097_ _1914_ _1916_ VGND VGND VPWR VPWR _2099_ sky130_fd_sc_hd__o211ai_4
X_5505_ _3631_ _2248_ _0950_ _0951_ VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__a22oi_1
X_6485_ _2011_ _2012_ _2022_ VGND VGND VPWR VPWR _2023_ sky130_fd_sc_hd__or3_4
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5436_ _0862_ _0875_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5367_ _0642_ _0768_ _0799_ _0800_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4318_ _3422_ VGND VGND VPWR VPWR _3423_ sky130_fd_sc_hd__clkbuf_4
X_5298_ _0205_ net38 _0596_ _0595_ _3718_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__a32oi_2
X_7106_ _2678_ _2697_ _2701_ VGND VGND VPWR VPWR _2702_ sky130_fd_sc_hd__nand3_1
X_4249_ _3352_ _3353_ _3354_ VGND VGND VPWR VPWR _3355_ sky130_fd_sc_hd__a21bo_1
X_7037_ _2457_ _2464_ VGND VGND VPWR VPWR _2627_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_383 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_843 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6270_ _1625_ _1754_ _1786_ VGND VGND VPWR VPWR _1787_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_121_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5221_ _0638_ _0639_ _0640_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__nand3_4
XFILLER_0_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5152_ _0296_ _0298_ _0422_ _0566_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4103_ _3210_ VGND VGND VPWR VPWR _3211_ sky130_fd_sc_hd__inv_2
X_5083_ net4 VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4034_ _0903_ _2051_ _3142_ VGND VGND VPWR VPWR _3143_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5985_ _1327_ _1474_ VGND VGND VPWR VPWR _1476_ sky130_fd_sc_hd__nor2_1
X_4936_ _0323_ _0329_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_75_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_10 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4867_ net178 net5 net6 _3242_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_21 _2412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_466 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6606_ _3196_ _3271_ _1854_ _1887_ VGND VGND VPWR VPWR _2155_ sky130_fd_sc_hd__and4_1
X_3818_ _0947_ VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4798_ _3723_ _0012_ _0179_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__a21o_1
X_6537_ _2074_ _2079_ VGND VGND VPWR VPWR _2080_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_7_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3749_ _0194_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__buf_4
XFILLER_0_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6468_ _2892_ _1898_ VGND VGND VPWR VPWR _2004_ sky130_fd_sc_hd__nand2_1
X_5419_ _0578_ _0839_ _0843_ _0857_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__a211oi_1
X_6399_ _1778_ _1797_ VGND VGND VPWR VPWR _1929_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5770_ _1232_ _1239_ _1240_ VGND VGND VPWR VPWR _1241_ sky130_fd_sc_hd__nand3_1
XFILLER_0_57_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4721_ _0019_ _0026_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__or2b_1
XFILLER_0_90_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4652_ _1264_ _0314_ net64 _3572_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__and4_1
XFILLER_0_71_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7440_ _2303_ _2309_ _3062_ _3064_ VGND VGND VPWR VPWR _3065_ sky130_fd_sc_hd__a31o_1
XFILLER_0_154_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput30 A[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_4
Xinput41 B[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_4
X_4583_ _2270_ _3685_ VGND VGND VPWR VPWR _3686_ sky130_fd_sc_hd__or2_1
X_7371_ _2974_ _2990_ VGND VGND VPWR VPWR _2992_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput52 B[27] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_2
XFILLER_0_4_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput63 B[8] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_2
XFILLER_0_12_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6322_ _1841_ _1842_ _1829_ VGND VGND VPWR VPWR _1845_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_776 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6253_ _1609_ _1610_ VGND VGND VPWR VPWR _1770_ sky130_fd_sc_hd__or2_1
X_5204_ _0614_ _0622_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__xnor2_2
X_6184_ _1686_ _1692_ _1693_ VGND VGND VPWR VPWR _1694_ sky130_fd_sc_hd__nand3_4
XFILLER_0_0_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5135_ _0321_ _0414_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__and2_1
X_5066_ _0346_ _0219_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4017_ _3108_ _3118_ VGND VGND VPWR VPWR _3126_ sky130_fd_sc_hd__nor2_2
XFILLER_0_137_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5968_ _1456_ _1305_ _1297_ VGND VGND VPWR VPWR _1457_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4919_ _3219_ _3220_ _3224_ _3225_ _3087_ _3486_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5899_ _1379_ _1380_ _1360_ _1361_ VGND VGND VPWR VPWR _1382_ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6940_ _2343_ _2349_ _2342_ VGND VGND VPWR VPWR _2520_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6871_ _2258_ _2261_ VGND VGND VPWR VPWR _2446_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5822_ _1942_ _1295_ VGND VGND VPWR VPWR _1298_ sky130_fd_sc_hd__nor2_1
X_5753_ _3430_ _2696_ _1219_ _1221_ VGND VGND VPWR VPWR _1223_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_57_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4704_ _0076_ _0077_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5684_ _0997_ _0895_ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7423_ _3136_ _3140_ _3138_ _3047_ _1723_ _1712_ VGND VGND VPWR VPWR _3048_ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4635_ _2675_ _3137_ _2237_ _2182_ _3046_ _3591_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__mux4_2
X_4566_ net139 _3667_ _3627_ VGND VGND VPWR VPWR _3669_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_114_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7354_ _2971_ _2972_ VGND VGND VPWR VPWR _2973_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6305_ _1651_ _1653_ _1824_ _1825_ VGND VGND VPWR VPWR _1826_ sky130_fd_sc_hd__o211ai_1
X_4497_ _3598_ _3599_ _3575_ VGND VGND VPWR VPWR _3601_ sky130_fd_sc_hd__a21oi_2
X_7285_ _3712_ _2880_ _3161_ VGND VGND VPWR VPWR _2897_ sky130_fd_sc_hd__o21ba_1
X_6236_ _1748_ _1749_ _1478_ VGND VGND VPWR VPWR _1751_ sky130_fd_sc_hd__o21a_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _1672_ _1673_ _1659_ VGND VGND VPWR VPWR _1675_ sky130_fd_sc_hd__a21o_1
X_5118_ _0526_ _0527_ net173 net202 VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__a211o_1
XFILLER_0_85_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6098_ _1597_ _1598_ VGND VGND VPWR VPWR _1600_ sky130_fd_sc_hd__nor2_1
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5049_ _0452_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_138_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_451 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4420_ _0085_ _1264_ _3195_ _3431_ VGND VGND VPWR VPWR _3524_ sky130_fd_sc_hd__nand4_1
XFILLER_0_53_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4351_ _3357_ _3359_ _3358_ VGND VGND VPWR VPWR _3456_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_50_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4282_ net31 net63 VGND VGND VPWR VPWR _3388_ sky130_fd_sc_hd__and2_4
XFILLER_0_10_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7070_ _2501_ _2662_ VGND VGND VPWR VPWR _2663_ sky130_fd_sc_hd__nor2_1
X_6021_ _1379_ _1381_ _1513_ _1514_ VGND VGND VPWR VPWR _1516_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_146_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6923_ _2443_ _2442_ VGND VGND VPWR VPWR _2502_ sky130_fd_sc_hd__and2b_1
XFILLER_0_49_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6854_ _2172_ _2174_ _2425_ _2426_ VGND VGND VPWR VPWR _2427_ sky130_fd_sc_hd__a211o_1
XFILLER_0_36_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3997_ _2335_ _2903_ VGND VGND VPWR VPWR _2914_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6785_ _2342_ _2343_ _2349_ VGND VGND VPWR VPWR _2351_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5805_ _0848_ _3200_ _3161_ VGND VGND VPWR VPWR _1280_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5736_ _3572_ _3651_ _2642_ _3422_ VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5667_ net136 _1127_ net119 net110 VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_32_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4618_ _3719_ VGND VGND VPWR VPWR _3720_ sky130_fd_sc_hd__clkbuf_4
X_7406_ _2346_ _1949_ VGND VGND VPWR VPWR _3030_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5598_ _1050_ _1051_ _1275_ net41 VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__and4bb_1
X_4549_ _3448_ _3537_ _3651_ _3449_ VGND VGND VPWR VPWR _3652_ sky130_fd_sc_hd__a22o_1
X_7337_ _2786_ _2792_ _2953_ VGND VGND VPWR VPWR _2954_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7268_ _3571_ _2702_ _2703_ _2867_ _2878_ VGND VGND VPWR VPWR _2879_ sky130_fd_sc_hd__a311o_1
X_6219_ _1720_ _1721_ _1731_ VGND VGND VPWR VPWR _1732_ sky130_fd_sc_hd__or3_4
X_7199_ _2643_ VGND VGND VPWR VPWR _2804_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3920_ _2040_ _2062_ _0936_ VGND VGND VPWR VPWR _2073_ sky130_fd_sc_hd__mux2_2
XFILLER_0_59_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3851_ _0303_ _0445_ VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3782_ _0554_ _0357_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6570_ _0861_ _3605_ VGND VGND VPWR VPWR _2116_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5521_ _0966_ _0967_ _0968_ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__nand3_1
XFILLER_0_26_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5452_ _0419_ _0879_ _0880_ _0889_ _0893_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__a311o_1
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4403_ _3305_ _3478_ _3479_ _3507_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__a31o_2
X_5383_ _0817_ _0818_ VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7122_ _2903_ _1767_ VGND VGND VPWR VPWR _2720_ sky130_fd_sc_hd__nand2_1
X_4334_ _3428_ _3438_ VGND VGND VPWR VPWR _3439_ sky130_fd_sc_hd__xor2_2
XFILLER_0_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7053_ _2624_ _2643_ _2644_ VGND VGND VPWR VPWR _2645_ sky130_fd_sc_hd__nor3_1
X_4265_ _3368_ _3369_ _3350_ VGND VGND VPWR VPWR _3371_ sky130_fd_sc_hd__o21a_1
X_6004_ _1495_ _1496_ VGND VGND VPWR VPWR _1497_ sky130_fd_sc_hd__xor2_2
X_4196_ _3156_ _3295_ _3302_ _3127_ VGND VGND VPWR VPWR _3303_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6906_ _2481_ _2482_ _2331_ _2332_ VGND VGND VPWR VPWR _2484_ sky130_fd_sc_hd__o211ai_2
X_6837_ _2171_ _2226_ _0721_ _0874_ VGND VGND VPWR VPWR _2408_ sky130_fd_sc_hd__nand4_1
XFILLER_0_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6768_ _2240_ _2267_ VGND VGND VPWR VPWR _2332_ sky130_fd_sc_hd__or2b_1
XFILLER_0_122_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5719_ _1054_ _1173_ _1183_ VGND VGND VPWR VPWR _1185_ sky130_fd_sc_hd__nand3_1
X_6699_ _1800_ _1977_ _2256_ VGND VGND VPWR VPWR _2257_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_646 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4050_ _2346_ _2903_ VGND VGND VPWR VPWR _3159_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput6 A[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4952_ _3442_ _3422_ _3511_ _2302_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__a22o_1
X_4883_ _0234_ _0235_ _0271_ _0272_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__or4bb_4
X_3903_ net14 VGND VGND VPWR VPWR _1887_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3834_ _0860_ _1122_ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6622_ _2718_ _0293_ _2170_ _2172_ VGND VGND VPWR VPWR _2173_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3765_ _0270_ _0368_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__or2_2
XFILLER_0_6_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6553_ _1914_ _1916_ _2096_ _2097_ VGND VGND VPWR VPWR _2098_ sky130_fd_sc_hd__a211o_1
XFILLER_0_144_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5504_ _3195_ _3633_ _2642_ _2686_ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__nand4_1
X_6484_ _2013_ _2021_ VGND VGND VPWR VPWR _2022_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5435_ _0874_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__buf_2
XFILLER_0_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5366_ _0797_ _0798_ _0778_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__a21oi_2
X_4317_ net64 VGND VGND VPWR VPWR _3422_ sky130_fd_sc_hd__buf_4
X_5297_ _0477_ _0688_ _0657_ _0656_ _0327_ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__a32o_1
X_7105_ net54 _2018_ VGND VGND VPWR VPWR _2701_ sky130_fd_sc_hd__or2b_1
X_4248_ net59 _0074_ net28 net58 VGND VGND VPWR VPWR _3354_ sky130_fd_sc_hd__a22o_1
X_7036_ _2453_ _2454_ _2466_ _2468_ VGND VGND VPWR VPWR _2626_ sky130_fd_sc_hd__a211o_1
X_4179_ _1209_ _3274_ _3204_ VGND VGND VPWR VPWR _3286_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_93_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5220_ _0506_ _0515_ _0514_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_11_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5151_ _3134_ _0337_ _0422_ _0564_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5082_ _0363_ _0364_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__nand2_1
X_4102_ _0903_ _3209_ VGND VGND VPWR VPWR _3210_ sky130_fd_sc_hd__or2b_2
X_4033_ _0903_ _2018_ VGND VGND VPWR VPWR _3142_ sky130_fd_sc_hd__and2b_1
XFILLER_0_154_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5984_ _1327_ _1474_ VGND VGND VPWR VPWR _1475_ sky130_fd_sc_hd__and2_2
XFILLER_0_136_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4935_ _1384_ _0328_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_11 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4866_ _0281_ _2642_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_22 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6605_ _1952_ _2001_ _2003_ _2004_ VGND VGND VPWR VPWR _2154_ sky130_fd_sc_hd__o2bb2a_1
X_3817_ _0936_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__clkbuf_4
X_4797_ _0178_ _3720_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3748_ net26 VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__clkbuf_4
X_6536_ _2077_ _2078_ VGND VGND VPWR VPWR _2079_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6467_ _1952_ _2001_ _2002_ VGND VGND VPWR VPWR _2003_ sky130_fd_sc_hd__a21bo_1
X_5418_ _0844_ _0847_ _0851_ _0853_ _0856_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__a311o_1
X_6398_ _1778_ _1797_ VGND VGND VPWR VPWR _1928_ sky130_fd_sc_hd__nor2_1
X_5349_ _3531_ net6 _0380_ _0161_ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7019_ _2564_ _2566_ _2605_ _2606_ VGND VGND VPWR VPWR _2607_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_97_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_814 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4720_ _0024_ _0025_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_674 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4651_ _0194_ _3422_ _3511_ _0324_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_83_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput20 A[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_4
XFILLER_0_72_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput31 A[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_25_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput64 B[9] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_4
X_4582_ _3620_ VGND VGND VPWR VPWR _3685_ sky130_fd_sc_hd__clkbuf_4
X_7370_ _2975_ _2989_ VGND VGND VPWR VPWR _2990_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput42 B[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput53 B[28] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_2
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6321_ _1829_ _1841_ _1842_ VGND VGND VPWR VPWR _1844_ sky130_fd_sc_hd__nand3_1
XFILLER_0_122_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_788 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6252_ _1761_ _1762_ _1765_ _1768_ VGND VGND VPWR VPWR _1769_ sky130_fd_sc_hd__or4_1
X_5203_ _0615_ _0621_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__xnor2_2
X_6183_ _1689_ _1691_ _1530_ _1532_ VGND VGND VPWR VPWR _1693_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_58_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5134_ _0321_ _0414_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5065_ _0469_ _0470_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__nor2_1
X_4016_ _1165_ _0630_ _1154_ _1144_ VGND VGND VPWR VPWR _3118_ sky130_fd_sc_hd__or4b_4
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5967_ _1297_ _1298_ VGND VGND VPWR VPWR _1456_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4918_ _3201_ _0196_ _0294_ _0307_ _0310_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__a221o_1
XFILLER_0_106_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5898_ _1360_ _1361_ _1379_ _1380_ VGND VGND VPWR VPWR _1381_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_145_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4849_ _0232_ _0233_ _0212_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6519_ _1034_ _1448_ _2057_ _2058_ VGND VGND VPWR VPWR _2060_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_608 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_663 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6870_ _2442_ _2443_ VGND VGND VPWR VPWR _2444_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5821_ _1942_ _1295_ VGND VGND VPWR VPWR _1297_ sky130_fd_sc_hd__and2_1
X_5752_ _1219_ _1221_ _3343_ _2686_ VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_17_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4703_ _3612_ _3675_ net151 VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_60_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5683_ net141 _0817_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7422_ _1067_ _1045_ _1034_ _1023_ _0914_ _0958_ VGND VGND VPWR VPWR _3047_ sky130_fd_sc_hd__mux4_1
X_4634_ _1111_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4565_ _3627_ _3666_ _3667_ VGND VGND VPWR VPWR _3668_ sky130_fd_sc_hd__and3_2
XFILLER_0_114_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7353_ _3591_ _2051_ VGND VGND VPWR VPWR _2972_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6304_ _2324_ net45 _1822_ _1823_ VGND VGND VPWR VPWR _1825_ sky130_fd_sc_hd__a22o_1
X_4496_ _3575_ _3598_ _3599_ VGND VGND VPWR VPWR _3600_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7284_ _1277_ _2880_ VGND VGND VPWR VPWR _2896_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6235_ _1478_ _1748_ _1749_ VGND VGND VPWR VPWR _1750_ sky130_fd_sc_hd__nor3_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _1659_ _1672_ _1673_ VGND VGND VPWR VPWR _1674_ sky130_fd_sc_hd__nand3_2
X_5117_ net173 net114 net125 _0527_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__o211ai_4
X_6097_ _1597_ _1598_ VGND VGND VPWR VPWR _1599_ sky130_fd_sc_hd__and2_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5048_ net40 VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__buf_2
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6999_ _2575_ _2583_ VGND VGND VPWR VPWR _2585_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4350_ _3450_ _3453_ _3447_ VGND VGND VPWR VPWR _3455_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4281_ _2127_ _3386_ VGND VGND VPWR VPWR _3387_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6020_ _1511_ _1512_ _1498_ VGND VGND VPWR VPWR _1514_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6922_ _2487_ VGND VGND VPWR VPWR _2501_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6853_ _2270_ _0688_ _2422_ _2424_ VGND VGND VPWR VPWR _2426_ sky130_fd_sc_hd__and4_1
XFILLER_0_49_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5804_ _3712_ _1270_ _1271_ _0309_ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_119_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6784_ _2342_ _2343_ _2349_ VGND VGND VPWR VPWR _2350_ sky130_fd_sc_hd__nand3_1
X_3996_ _2892_ VGND VGND VPWR VPWR _2903_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5735_ net64 _3572_ net3 _2642_ VGND VGND VPWR VPWR _1203_ sky130_fd_sc_hd__and4_1
XFILLER_0_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5666_ net119 net111 _1126_ _1127_ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__o211a_4
XFILLER_0_5_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4617_ _3718_ VGND VGND VPWR VPWR _3719_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7405_ _2829_ _2832_ VGND VGND VPWR VPWR _3029_ sky130_fd_sc_hd__or2b_1
XFILLER_0_44_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5597_ _1275_ _0654_ _1050_ _1051_ VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_5_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4548_ net3 VGND VGND VPWR VPWR _3651_ sky130_fd_sc_hd__clkbuf_4
X_7336_ _2787_ _2791_ VGND VGND VPWR VPWR _2953_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4479_ _3581_ _3582_ _3486_ VGND VGND VPWR VPWR _3583_ sky130_fd_sc_hd__mux2_1
X_7267_ _0844_ _2870_ _2873_ _2877_ VGND VGND VPWR VPWR _2878_ sky130_fd_sc_hd__a211o_1
X_6218_ _1722_ _1730_ VGND VGND VPWR VPWR _1731_ sky130_fd_sc_hd__xnor2_1
X_7198_ _2800_ _2801_ _2564_ _2704_ VGND VGND VPWR VPWR _2803_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_99_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6149_ _1653_ _1654_ VGND VGND VPWR VPWR _1655_ sky130_fd_sc_hd__nor2_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3850_ _1286_ _1296_ VGND VGND VPWR VPWR _1307_ sky130_fd_sc_hd__or2b_1
XFILLER_0_86_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3781_ _0303_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5520_ _0785_ _0786_ _0787_ VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_70_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5451_ _0890_ _0891_ _0575_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5382_ _0682_ net208 net140 VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__a21o_1
X_4402_ _2980_ _3484_ _3485_ _3506_ VGND VGND VPWR VPWR _3507_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7121_ _2716_ _2717_ VGND VGND VPWR VPWR _2719_ sky130_fd_sc_hd__nor2_1
X_4333_ _3429_ _3437_ VGND VGND VPWR VPWR _3438_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4264_ _3350_ _3368_ _3369_ VGND VGND VPWR VPWR _3370_ sky130_fd_sc_hd__nor3_2
XFILLER_0_1_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7052_ _2640_ _2641_ _2625_ _2626_ VGND VGND VPWR VPWR _2644_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6003_ _1330_ _1333_ VGND VGND VPWR VPWR _1496_ sky130_fd_sc_hd__or2_2
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4195_ _3296_ _3298_ _3299_ _3300_ _3077_ _3301_ VGND VGND VPWR VPWR _3302_ sky130_fd_sc_hd__mux4_1
XFILLER_0_66_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6905_ _2331_ _2332_ _2481_ _2482_ VGND VGND VPWR VPWR _2483_ sky130_fd_sc_hd__a211o_4
XFILLER_0_49_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6836_ _2226_ _0721_ _0874_ _2171_ VGND VGND VPWR VPWR _2407_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6767_ _2238_ _2239_ VGND VGND VPWR VPWR _2331_ sky130_fd_sc_hd__or2_1
X_3979_ _2707_ VGND VGND VPWR VPWR _2718_ sky130_fd_sc_hd__buf_4
X_5718_ _1054_ _1173_ _1183_ VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6698_ _1976_ _1970_ VGND VGND VPWR VPWR _2256_ sky130_fd_sc_hd__and2b_1
XFILLER_0_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5649_ _0390_ net11 _1854_ _0488_ VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_499 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7319_ _3133_ _0722_ VGND VGND VPWR VPWR _2934_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput7 A[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_2
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4951_ _2302_ _2368_ _3511_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__and3_1
X_4882_ _0268_ _0269_ _0148_ _0236_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_87_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3902_ _1865_ VGND VGND VPWR VPWR _1876_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6621_ _3720_ _0174_ _2762_ _2784_ VGND VGND VPWR VPWR _2172_ sky130_fd_sc_hd__nand4_2
X_3833_ _0870_ _1111_ VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3764_ _0303_ _0357_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6552_ _2093_ net182 _1988_ VGND VGND VPWR VPWR _2097_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5503_ _3431_ net4 net5 _3433_ VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__a22o_1
X_6483_ _2014_ _2020_ VGND VGND VPWR VPWR _2021_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_112_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5434_ _0873_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__buf_2
XFILLER_0_113_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5365_ _0778_ _0797_ _0798_ VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7104_ _2670_ _2698_ _2697_ VGND VGND VPWR VPWR _2700_ sky130_fd_sc_hd__o21ai_2
X_4316_ _3341_ _3349_ _3420_ VGND VGND VPWR VPWR _3421_ sky130_fd_sc_hd__o21ai_2
X_5296_ _1002_ _0722_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__nand2_2
XFILLER_0_11_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4247_ net59 _0074_ net28 VGND VGND VPWR VPWR _3353_ sky130_fd_sc_hd__and3_1
X_7035_ _2466_ VGND VGND VPWR VPWR _2625_ sky130_fd_sc_hd__inv_2
X_4178_ _3283_ _3284_ _1100_ VGND VGND VPWR VPWR _3285_ sky130_fd_sc_hd__mux2_2
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6819_ _2386_ _2387_ VGND VGND VPWR VPWR _2388_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_558 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5150_ _0328_ _3135_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__and2b_1
X_5081_ _0371_ _0392_ _0393_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__nand3_1
X_4101_ _1384_ VGND VGND VPWR VPWR _3209_ sky130_fd_sc_hd__clkbuf_8
X_4032_ _3132_ _3136_ _3138_ _3140_ _3077_ _1723_ VGND VGND VPWR VPWR _3141_ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5983_ _1335_ _1336_ VGND VGND VPWR VPWR _1474_ sky130_fd_sc_hd__and2b_1
XFILLER_0_74_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4934_ _0327_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_12 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4865_ _0249_ _0252_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_90_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3816_ _0521_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__clkbuf_4
X_6604_ _2015_ _2017_ VGND VGND VPWR VPWR _2153_ sky130_fd_sc_hd__or2_1
X_4796_ _2664_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3747_ _0172_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__clkbuf_4
X_6535_ _2160_ _0688_ _2075_ _2076_ VGND VGND VPWR VPWR _2078_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_803 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6466_ _0041_ net15 net16 _3645_ VGND VGND VPWR VPWR _2002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5417_ _0854_ _0826_ _0828_ _0855_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__a22o_1
X_6397_ _1787_ _1926_ VGND VGND VPWR VPWR _1927_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5348_ _0161_ _3531_ net6 VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__and3_1
X_5279_ _3589_ _0690_ _0000_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__o21bai_1
X_7018_ _2603_ _2604_ _2567_ _2568_ VGND VGND VPWR VPWR _2606_ sky130_fd_sc_hd__a211o_1
XFILLER_0_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4650_ _0477_ _3719_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput21 A[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_4
XFILLER_0_116_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput10 A[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_4
XFILLER_0_25_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput43 B[19] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
XFILLER_0_142_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput32 A[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_4
XFILLER_0_130_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput54 B[29] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_4
X_4581_ _3609_ net127 VGND VGND VPWR VPWR _3684_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6320_ _1838_ _1839_ _1840_ VGND VGND VPWR VPWR _1842_ sky130_fd_sc_hd__a21o_1
XFILLER_0_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput65 control[0] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6251_ _3414_ _1609_ _1610_ _0854_ _1766_ VGND VGND VPWR VPWR _1768_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5202_ _0618_ _0620_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__nor2_1
X_6182_ _1530_ _1532_ _1689_ _1691_ VGND VGND VPWR VPWR _1692_ sky130_fd_sc_hd__a211o_4
XFILLER_0_58_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_875 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5133_ _0544_ _0545_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5064_ _3440_ _0194_ _0339_ _0340_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__and4_1
XFILLER_0_79_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4015_ _0870_ VGND VGND VPWR VPWR _3108_ sky130_fd_sc_hd__buf_2
XFILLER_0_79_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5966_ _1454_ _1446_ _1303_ VGND VGND VPWR VPWR _1455_ sky130_fd_sc_hd__or3b_1
XFILLER_0_74_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4917_ _3712_ _0294_ _0295_ _0309_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__o22ai_1
X_5897_ _1363_ _1364_ _1378_ VGND VGND VPWR VPWR _1380_ sky130_fd_sc_hd__nor3_2
XFILLER_0_48_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4848_ _0212_ _0232_ _0233_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__nor3_1
XFILLER_0_75_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4779_ _0157_ _0158_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7498_ _3125_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__buf_6
X_6518_ _0226_ net48 _2057_ _2058_ VGND VGND VPWR VPWR _2059_ sky130_fd_sc_hd__nand4_1
XFILLER_0_43_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6449_ _1805_ _1981_ _1980_ VGND VGND VPWR VPWR _1983_ sky130_fd_sc_hd__a21o_1
XFILLER_0_100_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5820_ _1294_ VGND VGND VPWR VPWR _1295_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5751_ _3633_ net6 _0380_ _3195_ VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_127_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4702_ _0073_ _0075_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5682_ _0549_ net164 _0553_ _1145_ VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__a31o_1
XFILLER_0_72_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7421_ _2886_ _3045_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__nand2_2
XFILLER_0_154_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_678 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4633_ _3490_ _3486_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4564_ _3664_ _3665_ _3548_ net155 VGND VGND VPWR VPWR _3667_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_103_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7352_ _3490_ _2018_ VGND VGND VPWR VPWR _2971_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7283_ _0309_ _2882_ _2883_ _3589_ VGND VGND VPWR VPWR _2895_ sky130_fd_sc_hd__o22a_1
X_6303_ _2324_ _1007_ _1822_ _1823_ VGND VGND VPWR VPWR _1824_ sky130_fd_sc_hd__nand4_2
X_4495_ _3395_ _3396_ _3482_ _3389_ VGND VGND VPWR VPWR _3599_ sky130_fd_sc_hd__a211o_1
XFILLER_0_12_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6234_ _1746_ _1747_ _1586_ _1588_ VGND VGND VPWR VPWR _1749_ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _1669_ _1670_ _1671_ VGND VGND VPWR VPWR _1673_ sky130_fd_sc_hd__a21o_1
X_5116_ _0486_ _0487_ _0524_ _0525_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__a2bb2o_1
X_6096_ _1435_ _1434_ VGND VGND VPWR VPWR _1598_ sky130_fd_sc_hd__or2_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5047_ _0341_ _0343_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__or2_1
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6998_ _2575_ _2583_ VGND VGND VPWR VPWR _2584_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5949_ _1434_ _1436_ VGND VGND VPWR VPWR _1437_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4280_ _3385_ VGND VGND VPWR VPWR _3386_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6921_ _2326_ _2490_ VGND VGND VPWR VPWR _2500_ sky130_fd_sc_hd__nand2_1
X_6852_ _2270_ _0689_ _2422_ _2424_ VGND VGND VPWR VPWR _2425_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_49_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5803_ _0438_ _1271_ _1277_ VGND VGND VPWR VPWR _1278_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6783_ _2347_ _2348_ VGND VGND VPWR VPWR _2349_ sky130_fd_sc_hd__xnor2_1
X_3995_ _2881_ VGND VGND VPWR VPWR _2892_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5734_ _1200_ _1201_ VGND VGND VPWR VPWR _1202_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5665_ _1088_ _1090_ _1124_ _1125_ VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4616_ net36 VGND VGND VPWR VPWR _3718_ sky130_fd_sc_hd__buf_2
XFILLER_0_5_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7404_ _3026_ _3027_ VGND VGND VPWR VPWR _3028_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_143_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5596_ _0085_ _2302_ _0325_ _0452_ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__and4_1
X_7335_ _2766_ _2799_ _2765_ VGND VGND VPWR VPWR _2952_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_5_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4547_ _0292_ net32 VGND VGND VPWR VPWR _3650_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4478_ _3219_ _3225_ _1100_ VGND VGND VPWR VPWR _3582_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7266_ _0575_ _2874_ _2875_ _2876_ VGND VGND VPWR VPWR _2877_ sky130_fd_sc_hd__a211o_1
XFILLER_0_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6217_ _1724_ _1729_ VGND VGND VPWR VPWR _1730_ sky130_fd_sc_hd__xnor2_1
X_7197_ _2564_ _2704_ _2800_ _2801_ VGND VGND VPWR VPWR _2802_ sky130_fd_sc_hd__o211a_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ _0106_ _1007_ _1651_ _1652_ VGND VGND VPWR VPWR _1654_ sky130_fd_sc_hd__o2bb2a_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ _1541_ _1542_ _1577_ _1578_ VGND VGND VPWR VPWR _1579_ sky130_fd_sc_hd__or4bb_4
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsplit70 _0074_ VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__buf_6
X_3780_ _0455_ _0510_ _0532_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5450_ _0848_ _0884_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4401_ _3489_ _3495_ _3499_ _3505_ VGND VGND VPWR VPWR _3506_ sky130_fd_sc_hd__or4b_1
XFILLER_0_2_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5381_ _0814_ _0815_ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__nor2b_1
XFILLER_0_10_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7120_ _0172_ _0052_ _1799_ net20 VGND VGND VPWR VPWR _2717_ sky130_fd_sc_hd__and4_1
X_4332_ _3435_ _3436_ VGND VGND VPWR VPWR _3437_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4263_ _3365_ _3366_ _3367_ VGND VGND VPWR VPWR _3369_ sky130_fd_sc_hd__a21oi_1
X_7051_ _2625_ _2626_ _2640_ _2641_ VGND VGND VPWR VPWR _2643_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_66_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6002_ _1491_ _1494_ VGND VGND VPWR VPWR _1495_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4194_ _1723_ VGND VGND VPWR VPWR _3301_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6904_ _2479_ _2480_ _2444_ VGND VGND VPWR VPWR _2482_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6835_ _2404_ _2405_ VGND VGND VPWR VPWR _2406_ sky130_fd_sc_hd__or2_1
XFILLER_0_135_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_559 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3978_ _2696_ VGND VGND VPWR VPWR _2707_ sky130_fd_sc_hd__buf_4
XFILLER_0_58_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6766_ _1982_ _2266_ VGND VGND VPWR VPWR _2330_ sky130_fd_sc_hd__and2b_1
X_5717_ _1174_ _1182_ VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__xnor2_1
X_6697_ _2243_ _2254_ VGND VGND VPWR VPWR _2255_ sky130_fd_sc_hd__xor2_1
XFILLER_0_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5648_ _3451_ _3452_ _2598_ _1854_ VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__nand4_2
XFILLER_0_5_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5579_ _1026_ _1031_ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7318_ _2675_ _0875_ VGND VGND VPWR VPWR _2933_ sky130_fd_sc_hd__nand2_1
X_7249_ _2857_ _2858_ VGND VGND VPWR VPWR _2859_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput8 A[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_127_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_523 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4950_ _0095_ _0110_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4881_ _0148_ _0236_ _0268_ _0269_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__a211o_1
X_3901_ _1854_ VGND VGND VPWR VPWR _1865_ sky130_fd_sc_hd__buf_4
XFILLER_0_145_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6620_ _0174_ _2751_ _2784_ _3719_ VGND VGND VPWR VPWR _2170_ sky130_fd_sc_hd__a22o_1
X_3832_ _0925_ _0969_ _1012_ _1089_ _1100_ VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__o32a_1
XFILLER_0_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6551_ _1988_ _2093_ _2094_ VGND VGND VPWR VPWR _2096_ sky130_fd_sc_hd__and3_1
XFILLER_0_144_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5502_ _2892_ _2707_ _0781_ _0780_ _2773_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__a32o_1
XFILLER_0_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3763_ _0346_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__buf_4
X_6482_ _2017_ _2019_ VGND VGND VPWR VPWR _2020_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5433_ net43 VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__buf_2
XFILLER_0_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5364_ _0793_ _0795_ _0796_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4315_ _3348_ _3342_ VGND VGND VPWR VPWR _3420_ sky130_fd_sc_hd__or2b_1
XFILLER_0_11_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7103_ _2670_ _2697_ _2698_ VGND VGND VPWR VPWR _2699_ sky130_fd_sc_hd__or3_1
X_5295_ _0721_ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__clkbuf_4
X_4246_ net58 VGND VGND VPWR VPWR _3352_ sky130_fd_sc_hd__clkbuf_4
X_7034_ _2622_ _2623_ VGND VGND VPWR VPWR _2624_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4177_ _1034_ _1045_ _1067_ _3209_ _0914_ _0958_ VGND VGND VPWR VPWR _3284_ sky130_fd_sc_hd__mux4_2
XFILLER_0_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6818_ _3685_ _2510_ _2177_ _2176_ VGND VGND VPWR VPWR _2387_ sky130_fd_sc_hd__a31o_1
XFILLER_0_65_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6749_ _2303_ _2309_ VGND VGND VPWR VPWR _2311_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_618 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5080_ _0484_ _0485_ _0465_ _0467_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__o211a_1
X_4100_ _1045_ _1067_ _0914_ VGND VGND VPWR VPWR _3208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4031_ _2346_ _2412_ _3139_ _2138_ _0914_ _0958_ VGND VGND VPWR VPWR _3140_ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5982_ _1320_ _1322_ VGND VGND VPWR VPWR _1473_ sky130_fd_sc_hd__nor2_2
XFILLER_0_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4933_ _0326_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__buf_2
XFILLER_0_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4864_ _0250_ _0251_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__nor2_1
XANTENNA_13 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6603_ net152 _2148_ _2150_ VGND VGND VPWR VPWR _2152_ sky130_fd_sc_hd__a21oi_2
X_4795_ _0175_ _0176_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__nand2_1
X_3815_ _0914_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3746_ _0161_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__buf_6
XFILLER_0_70_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6534_ _2075_ _2076_ _2160_ _0688_ VGND VGND VPWR VPWR _2077_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6465_ _3645_ _0041_ net15 VGND VGND VPWR VPWR _2001_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_815 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5416_ _3414_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6396_ _1789_ _1925_ VGND VGND VPWR VPWR _1926_ sky130_fd_sc_hd__xor2_1
XFILLER_0_100_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5347_ _0042_ _2696_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5278_ _3128_ _0689_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__or2_1
X_4229_ net192 _3335_ VGND VGND VPWR VPWR _3336_ sky130_fd_sc_hd__xor2_1
X_7017_ _2567_ _2568_ _2603_ _2604_ VGND VGND VPWR VPWR _2605_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_98_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4580_ _3609_ net126 VGND VGND VPWR VPWR _3683_ sky130_fd_sc_hd__or2_1
Xinput11 A[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_25_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput22 A[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_4
Xinput44 B[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_6
Xinput55 B[2] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_142_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput33 B[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_8
Xinput66 control[1] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_2
XFILLER_0_80_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6250_ _0199_ _3727_ _3487_ _3161_ VGND VGND VPWR VPWR _1766_ sky130_fd_sc_hd__o31a_1
XFILLER_0_110_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5201_ _3631_ _0247_ _0616_ _0617_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__o2bb2a_1
X_6181_ _3620_ _2707_ _1687_ _1688_ VGND VGND VPWR VPWR _1691_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_58_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5132_ _0540_ _0541_ _0542_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5063_ _3440_ _0339_ _0099_ _1275_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_79_415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4014_ _3035_ _3056_ _3066_ _3087_ VGND VGND VPWR VPWR _3097_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_74_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5965_ _1450_ _1451_ VGND VGND VPWR VPWR _1454_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4916_ _0308_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__clkbuf_4
X_5896_ _1363_ _1364_ _1378_ VGND VGND VPWR VPWR _1379_ sky130_fd_sc_hd__o21a_2
X_4847_ _0213_ _0214_ _0231_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__nor3_1
XFILLER_0_90_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4778_ net116 _0156_ _0093_ _0067_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7497_ net92 _2886_ _3045_ _3124_ VGND VGND VPWR VPWR _3125_ sky130_fd_sc_hd__and4b_2
XFILLER_0_43_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6517_ _2324_ _1169_ _1295_ _0106_ VGND VGND VPWR VPWR _2058_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6448_ _1805_ _1980_ _1981_ VGND VGND VPWR VPWR _1982_ sky130_fd_sc_hd__nand3_2
XFILLER_0_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6379_ _1884_ _1885_ _1905_ _1906_ VGND VGND VPWR VPWR _1907_ sky130_fd_sc_hd__or4_4
XFILLER_0_101_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5750_ _3433_ _3270_ net6 net7 VGND VGND VPWR VPWR _1219_ sky130_fd_sc_hd__and4_1
XFILLER_0_57_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4701_ _0071_ _0072_ net212 _3672_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__a211o_1
X_5681_ _0821_ _1143_ VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__or2_4
XFILLER_0_84_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4632_ _3589_ _3722_ _0000_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7420_ _0181_ _2888_ _2889_ _2899_ _3044_ VGND VGND VPWR VPWR _3045_ sky130_fd_sc_hd__o311a_1
XFILLER_0_44_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4563_ _3548_ _3628_ _3664_ _3665_ VGND VGND VPWR VPWR _3666_ sky130_fd_sc_hd__a211o_1
XFILLER_0_80_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7351_ _2956_ _2968_ VGND VGND VPWR VPWR _2970_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4494_ _3480_ _3597_ VGND VGND VPWR VPWR _3598_ sky130_fd_sc_hd__nor2_1
X_6302_ _3530_ _0720_ _0873_ _2379_ VGND VGND VPWR VPWR _1823_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7282_ _0844_ _2893_ VGND VGND VPWR VPWR _2894_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6233_ _1586_ _1588_ _1746_ _1747_ VGND VGND VPWR VPWR _1748_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _1669_ _1670_ _1671_ VGND VGND VPWR VPWR _1672_ sky130_fd_sc_hd__nand3_1
X_5115_ _0486_ _0487_ _0524_ _0525_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__or4bb_4
X_6095_ _1594_ _1596_ VGND VGND VPWR VPWR _1597_ sky130_fd_sc_hd__xnor2_4
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5046_ _1384_ _0328_ _0323_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6997_ _2581_ _2582_ VGND VGND VPWR VPWR _2583_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5948_ _1138_ _1265_ _1435_ VGND VGND VPWR VPWR _1436_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5879_ _1207_ _1210_ VGND VGND VPWR VPWR _1360_ sky130_fd_sc_hd__or2b_1
XFILLER_0_36_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_690 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6920_ _0419_ _2307_ _2325_ _2498_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__a211o_4
XFILLER_0_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6851_ _2664_ _2718_ _0328_ _0454_ VGND VGND VPWR VPWR _2424_ sky130_fd_sc_hd__nand4_1
XFILLER_0_49_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5802_ _0000_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__clkbuf_4
X_3994_ net60 VGND VGND VPWR VPWR _2881_ sky130_fd_sc_hd__clkbuf_4
X_6782_ _2903_ _1952_ VGND VGND VPWR VPWR _2348_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5733_ _2445_ _0220_ _1197_ _1199_ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5664_ net118 _1090_ _1124_ _1125_ VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4615_ _3305_ _3683_ _3684_ _3717_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__a31o_2
XFILLER_0_60_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5595_ _3635_ _0325_ _0452_ _3440_ VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_5_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7403_ _2779_ _2780_ _2782_ VGND VGND VPWR VPWR _3027_ sky130_fd_sc_hd__a21oi_1
X_4546_ _3643_ _3648_ VGND VGND VPWR VPWR _3649_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7334_ _3134_ _0559_ _0420_ _2950_ VGND VGND VPWR VPWR _2951_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4477_ _3220_ _3221_ _3077_ VGND VGND VPWR VPWR _3581_ sky130_fd_sc_hd__mux2_1
X_7265_ _0855_ _2694_ _2695_ _0854_ VGND VGND VPWR VPWR _2876_ sky130_fd_sc_hd__a22o_1
X_6216_ _1727_ _1728_ VGND VGND VPWR VPWR _1729_ sky130_fd_sc_hd__or2_1
X_7196_ _2765_ _2766_ _2799_ VGND VGND VPWR VPWR _2801_ sky130_fd_sc_hd__a21o_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6147_ _1651_ _1652_ _0106_ net45 VGND VGND VPWR VPWR _1653_ sky130_fd_sc_hd__and4bb_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ _1575_ _1576_ _1413_ _1543_ VGND VGND VPWR VPWR _1578_ sky130_fd_sc_hd__a211o_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5029_ _0428_ _0430_ _0431_ _3587_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__o211a_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4400_ _0860_ _3503_ _3504_ _3481_ VGND VGND VPWR VPWR _3505_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5380_ _0812_ _0813_ _0673_ _0718_ VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__a211o_1
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4331_ net163 _3343_ _3432_ _3434_ VGND VGND VPWR VPWR _3436_ sky130_fd_sc_hd__and4_1
XFILLER_0_67_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4262_ _3365_ _3366_ _3367_ VGND VGND VPWR VPWR _3368_ sky130_fd_sc_hd__and3_4
XFILLER_0_10_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7050_ _2638_ _2639_ _2462_ _2627_ VGND VGND VPWR VPWR _2641_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6001_ _0215_ _1007_ _1492_ _1490_ VGND VGND VPWR VPWR _1494_ sky130_fd_sc_hd__a22oi_1
X_4193_ _3139_ _2138_ _2182_ _2237_ _0903_ _0958_ VGND VGND VPWR VPWR _3300_ sky130_fd_sc_hd__mux4_1
XFILLER_0_66_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6903_ _2444_ _2479_ _2480_ VGND VGND VPWR VPWR _2481_ sky130_fd_sc_hd__and3_2
XFILLER_0_148_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6834_ _2402_ _1448_ _2335_ _2400_ VGND VGND VPWR VPWR _2405_ sky130_fd_sc_hd__and4b_1
XFILLER_0_119_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3977_ _2686_ VGND VGND VPWR VPWR _2696_ sky130_fd_sc_hd__buf_6
XFILLER_0_58_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6765_ _2265_ _2241_ VGND VGND VPWR VPWR _2329_ sky130_fd_sc_hd__and2b_1
XFILLER_0_135_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5716_ _1180_ _1181_ VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6696_ _2244_ _2253_ VGND VGND VPWR VPWR _2254_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_143_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5647_ _0281_ net10 VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5578_ _0419_ _1028_ _1029_ _1030_ _0575_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__a32o_1
XFILLER_0_130_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4529_ net61 VGND VGND VPWR VPWR _3632_ sky130_fd_sc_hd__buf_4
X_7317_ _0174_ _2587_ VGND VGND VPWR VPWR _2932_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7248_ _2654_ _2657_ _2856_ VGND VGND VPWR VPWR _2858_ sky130_fd_sc_hd__or3_1
X_7179_ _2774_ _2781_ VGND VGND VPWR VPWR _2782_ sky130_fd_sc_hd__nor2_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput9 A[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_2
XFILLER_0_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4880_ _0266_ _0267_ _0246_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__a21oi_1
X_3900_ net13 VGND VGND VPWR VPWR _1854_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3831_ _0980_ VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6550_ _2091_ _2092_ _1910_ _1989_ VGND VGND VPWR VPWR _2094_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3762_ _0335_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5501_ _0773_ _0774_ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6481_ _3385_ _2576_ _2015_ _2016_ VGND VGND VPWR VPWR _2019_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_70_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_777 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5432_ _0861_ _0868_ _0871_ _0844_ VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__o211a_1
X_5363_ _0793_ _0795_ _0796_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__nand3_4
XFILLER_0_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4314_ _3340_ _3372_ _3373_ VGND VGND VPWR VPWR _3419_ sky130_fd_sc_hd__nor3_1
XFILLER_0_11_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7102_ _2681_ _2673_ VGND VGND VPWR VPWR _2698_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5294_ _0720_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__buf_2
X_4245_ _0194_ net60 VGND VGND VPWR VPWR _3351_ sky130_fd_sc_hd__nand2_1
X_7033_ _2614_ _2621_ VGND VGND VPWR VPWR _2623_ sky130_fd_sc_hd__and2_1
X_4176_ _3139_ _2412_ _2346_ _1023_ _0925_ _0969_ VGND VGND VPWR VPWR _3283_ sky130_fd_sc_hd__mux4_2
XFILLER_0_117_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6817_ _2384_ _2385_ VGND VGND VPWR VPWR _2386_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_618 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6748_ _2303_ _2309_ VGND VGND VPWR VPWR _2310_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6679_ _2191_ _2192_ _2233_ _2234_ VGND VGND VPWR VPWR _2235_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_116_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4030_ _2456_ VGND VGND VPWR VPWR _3139_ sky130_fd_sc_hd__buf_4
XFILLER_0_154_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5981_ _0861_ _1461_ _1465_ _1470_ VGND VGND VPWR VPWR _1472_ sky130_fd_sc_hd__a211o_1
XFILLER_0_149_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_803 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4932_ _0325_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4863_ _0161_ _3531_ _3537_ _3651_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__and4_1
X_6602_ _2147_ _2148_ _2150_ VGND VGND VPWR VPWR _2151_ sky130_fd_sc_hd__and3_2
XANTENNA_14 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3814_ _0903_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__buf_4
X_4794_ _2718_ _0174_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3745_ net58 VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__buf_8
X_6533_ _2259_ _0327_ _0454_ _2226_ VGND VGND VPWR VPWR _2076_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6464_ _1995_ _1997_ _1998_ VGND VGND VPWR VPWR _2000_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5415_ _3194_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6395_ _1923_ _1924_ VGND VGND VPWR VPWR _1925_ sky130_fd_sc_hd__xor2_4
XFILLER_0_112_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5346_ _0769_ _0777_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__xor2_2
XFILLER_0_11_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5277_ _1723_ _0701_ _0702_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4228_ net145 _3259_ VGND VGND VPWR VPWR _3335_ sky130_fd_sc_hd__nand2_1
X_7016_ _2601_ _2602_ _2569_ _2393_ VGND VGND VPWR VPWR _2604_ sky130_fd_sc_hd__o211ai_4
X_4159_ _3215_ _3264_ _3266_ VGND VGND VPWR VPWR _3267_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput12 A[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_6
XFILLER_0_24_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput34 B[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_142_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput23 A[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_6
Xinput45 B[20] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput56 B[30] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_8
Xinput67 control[2] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_4
XFILLER_0_52_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5200_ _0616_ _0617_ _3631_ _0247_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__and4bb_1
X_6180_ _3619_ _2696_ _1687_ _1688_ VGND VGND VPWR VPWR _1689_ sky130_fd_sc_hd__and4_2
X_5131_ _0540_ _0541_ _0542_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5062_ _0360_ _0367_ _0366_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__a21bo_1
X_4013_ _3077_ VGND VGND VPWR VPWR _3087_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5964_ _1303_ _1447_ _1452_ VGND VGND VPWR VPWR _1453_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4915_ net65 _1144_ _1154_ _1165_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__or4b_1
X_5895_ _1369_ _1377_ VGND VGND VPWR VPWR _1378_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4846_ _0213_ _0214_ _0231_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4777_ _0093_ _0067_ net116 _0156_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_105_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6516_ _0117_ _2335_ _1170_ _1295_ VGND VGND VPWR VPWR _2057_ sky130_fd_sc_hd__nand4_2
X_7496_ net84 _3112_ _3122_ _3123_ VGND VGND VPWR VPWR _3124_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6447_ _1631_ _1807_ VGND VGND VPWR VPWR _1981_ sky130_fd_sc_hd__or2_1
X_6378_ _1903_ _1904_ _1692_ _1694_ VGND VGND VPWR VPWR _1906_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5329_ _0755_ _0758_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_100_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4700_ net212 _3672_ _0071_ _0072_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__o211ai_4
X_5680_ _0819_ _0997_ VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__or2b_1
XFILLER_0_84_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4631_ _3204_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__buf_2
XFILLER_0_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4562_ _3662_ _3663_ _3642_ VGND VGND VPWR VPWR _3665_ sky130_fd_sc_hd__a21oi_2
X_7350_ _2964_ _2967_ VGND VGND VPWR VPWR _2968_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4493_ _2182_ _3425_ _2138_ _3386_ VGND VGND VPWR VPWR _3597_ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7281_ _3285_ _0435_ _1467_ _2891_ _0867_ _0573_ VGND VGND VPWR VPWR _2893_ sky130_fd_sc_hd__mux4_1
X_6301_ _2379_ _2445_ _0720_ _0873_ VGND VGND VPWR VPWR _1822_ sky130_fd_sc_hd__nand4_2
X_6232_ _1743_ _1744_ _1641_ VGND VGND VPWR VPWR _1747_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6163_ _1500_ _1508_ _1507_ VGND VGND VPWR VPWR _1671_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _0522_ _0523_ _0392_ _0489_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__o211ai_2
X_6094_ _1319_ _1433_ _1595_ VGND VGND VPWR VPWR _1596_ sky130_fd_sc_hd__a21oi_4
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _0354_ _0356_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6996_ _2171_ _2226_ _0722_ _0875_ _2410_ VGND VGND VPWR VPWR _2582_ sky130_fd_sc_hd__a41o_1
XFILLER_0_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5947_ _1262_ _1263_ VGND VGND VPWR VPWR _1435_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5878_ _1215_ _1216_ _1249_ _1250_ VGND VGND VPWR VPWR _1359_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_145_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4829_ _0123_ _0127_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__and2b_1
XFILLER_0_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7479_ _1592_ _1603_ _1668_ VGND VGND VPWR VPWR _3106_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6850_ _2707_ _0327_ _0454_ _2664_ VGND VGND VPWR VPWR _2422_ sky130_fd_sc_hd__a22o_1
X_6781_ _2344_ _2345_ VGND VGND VPWR VPWR _2347_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5801_ _1272_ _1274_ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__xor2_1
XFILLER_0_9_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3993_ _0619_ _0652_ _0663_ _2861_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__a31o_1
XFILLER_0_85_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5732_ _3530_ net38 _1197_ _1199_ VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__nand4_2
XFILLER_0_45_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5663_ _1121_ _1123_ _0975_ _1091_ VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_72_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4614_ _0652_ _3691_ _3693_ _3716_ VGND VGND VPWR VPWR _3717_ sky130_fd_sc_hd__a31o_1
XFILLER_0_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5594_ _0908_ _0910_ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7402_ _1067_ net54 _2809_ _2808_ VGND VGND VPWR VPWR _3026_ sky130_fd_sc_hd__a31o_1
XFILLER_0_143_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4545_ _3646_ _3647_ VGND VGND VPWR VPWR _3648_ sky130_fd_sc_hd__nor2_1
X_7333_ _3133_ _0689_ _2789_ VGND VGND VPWR VPWR _2950_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap120 _1904_ VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__buf_1
XFILLER_0_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4476_ _3127_ VGND VGND VPWR VPWR _3580_ sky130_fd_sc_hd__buf_2
X_7264_ _0313_ _2319_ VGND VGND VPWR VPWR _2875_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6215_ _3430_ _2499_ _1725_ _1726_ VGND VGND VPWR VPWR _1728_ sky130_fd_sc_hd__o2bb2a_1
X_7195_ _2765_ _2766_ _2799_ VGND VGND VPWR VPWR _2800_ sky130_fd_sc_hd__nand3_1
XFILLER_0_0_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6146_ _2379_ _0720_ _0873_ _2313_ VGND VGND VPWR VPWR _1652_ sky130_fd_sc_hd__a22oi_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6077_ _1413_ net121 _1575_ _1576_ VGND VGND VPWR VPWR _1577_ sky130_fd_sc_hd__o211ai_4
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5028_ _3144_ _0196_ _3727_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__o21ai_1
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6979_ _2536_ _2537_ _2560_ _2561_ VGND VGND VPWR VPWR _2563_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_614 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4330_ _0423_ _3430_ _3432_ _3434_ VGND VGND VPWR VPWR _3435_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_50_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4261_ _3315_ _3323_ _3322_ VGND VGND VPWR VPWR _3367_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_10_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6000_ _1489_ VGND VGND VPWR VPWR _1492_ sky130_fd_sc_hd__inv_2
X_4192_ _3137_ _2675_ _3133_ _2762_ _0903_ _0958_ VGND VGND VPWR VPWR _3299_ sky130_fd_sc_hd__mux4_1
XFILLER_0_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6902_ _2476_ _2477_ _2446_ _2447_ VGND VGND VPWR VPWR _2480_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_49_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6833_ _2335_ _1448_ _2400_ _2403_ VGND VGND VPWR VPWR _2404_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3976_ net5 VGND VGND VPWR VPWR _2686_ sky130_fd_sc_hd__buf_4
XFILLER_0_64_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6764_ _2131_ _2272_ VGND VGND VPWR VPWR _2328_ sky130_fd_sc_hd__and2b_1
XFILLER_0_116_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5715_ _1178_ _1179_ _1074_ _1076_ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_18_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6695_ _2245_ _2252_ VGND VGND VPWR VPWR _2253_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_143_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5646_ _1104_ _1105_ VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__xor2_1
XFILLER_0_61_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_466 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5577_ _0573_ _2095_ _0890_ VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4528_ _3343_ VGND VGND VPWR VPWR _3631_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7316_ _3139_ _1448_ _2771_ _2770_ VGND VGND VPWR VPWR _2931_ sky130_fd_sc_hd__a31o_1
X_4459_ _3379_ _3472_ VGND VGND VPWR VPWR _3563_ sky130_fd_sc_hd__or2_1
X_7247_ _2654_ _2657_ _2856_ VGND VGND VPWR VPWR _2857_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7178_ _2779_ _2780_ VGND VGND VPWR VPWR _2781_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6129_ _1631_ _1632_ VGND VGND VPWR VPWR _1633_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3830_ _1078_ VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__inv_2
X_3761_ _0324_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5500_ _0778_ _0797_ _0798_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__nand3_2
XFILLER_0_55_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6480_ _2015_ _2016_ _3385_ _2576_ VGND VGND VPWR VPWR _2017_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_54_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5431_ _0848_ _0869_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5362_ _0628_ _0637_ _0636_ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_140_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4313_ _3305_ _3383_ _3384_ _3418_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__a31o_2
XFILLER_0_10_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7101_ _2694_ _2695_ VGND VGND VPWR VPWR _2697_ sky130_fd_sc_hd__nor2_2
X_5293_ net42 VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__buf_2
XFILLER_0_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7032_ _2614_ _2621_ VGND VGND VPWR VPWR _2622_ sky130_fd_sc_hd__nor2_1
X_4244_ _3341_ _3349_ VGND VGND VPWR VPWR _3350_ sky130_fd_sc_hd__xnor2_2
X_4175_ _3276_ _3281_ VGND VGND VPWR VPWR _3282_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6816_ _3685_ _2543_ VGND VGND VPWR VPWR _2385_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6747_ _2280_ _2296_ _2308_ VGND VGND VPWR VPWR _2309_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3959_ _2489_ VGND VGND VPWR VPWR _2499_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6678_ _2231_ _2232_ _2194_ _2195_ VGND VGND VPWR VPWR _2234_ sky130_fd_sc_hd__a211o_1
XFILLER_0_104_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5629_ _1071_ _1072_ _1085_ VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__nor3_2
XFILLER_0_61_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5980_ _3295_ _1469_ _0861_ VGND VGND VPWR VPWR _1470_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4931_ net39 VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__clkbuf_4
X_4862_ _3531_ _3537_ _2248_ _3645_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_75_815 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_528 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6601_ _2000_ _2005_ _1999_ VGND VGND VPWR VPWR _2150_ sky130_fd_sc_hd__a21bo_1
X_3813_ _0892_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4793_ _3133_ _0174_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_15 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3744_ _0128_ _0139_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__or2_1
X_6532_ _2215_ _2259_ _0327_ _0454_ VGND VGND VPWR VPWR _2075_ sky130_fd_sc_hd__and4_1
X_6463_ _1995_ _1997_ _1998_ VGND VGND VPWR VPWR _1999_ sky130_fd_sc_hd__nand3_1
XFILLER_0_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput100 net100 VGND VGND VPWR VPWR result[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5414_ _0828_ _0852_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6394_ _1748_ _1750_ VGND VGND VPWR VPWR _1924_ sky130_fd_sc_hd__nor2_2
XFILLER_0_100_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5345_ _0770_ _0776_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_56_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5276_ _1100_ _3145_ _3492_ _1723_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4227_ net193 _3333_ VGND VGND VPWR VPWR _3334_ sky130_fd_sc_hd__xnor2_2
X_7015_ _2569_ _2393_ _2601_ _2602_ VGND VGND VPWR VPWR _2603_ sky130_fd_sc_hd__a211o_2
X_4158_ _3215_ _3264_ _3265_ VGND VGND VPWR VPWR _3266_ sky130_fd_sc_hd__a21oi_1
X_4089_ _3196_ VGND VGND VPWR VPWR _3197_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_829 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput13 A[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_4
XFILLER_0_141_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput46 B[21] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_4
Xinput24 A[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput35 B[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_2
XFILLER_0_141_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput68 control[3] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_2
XFILLER_0_52_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput57 B[31] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5130_ _0283_ _0282_ _0410_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__nor3_1
X_5061_ _0344_ _0352_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__or2b_1
X_4012_ _1712_ VGND VGND VPWR VPWR _3077_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5963_ _1450_ _1451_ VGND VGND VPWR VPWR _1452_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4914_ net124 _0295_ _3204_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5894_ _1375_ _1376_ VGND VGND VPWR VPWR _1377_ sky130_fd_sc_hd__xor2_2
XFILLER_0_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4845_ _0222_ _0230_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4776_ _0119_ _0120_ _0153_ _0154_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6515_ _1841_ _1844_ VGND VGND VPWR VPWR _2056_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7495_ net88 _2669_ _2676_ _2692_ VGND VGND VPWR VPWR _3123_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_141_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6446_ _1802_ _1979_ VGND VGND VPWR VPWR _1980_ sky130_fd_sc_hd__xor2_1
XFILLER_0_101_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6377_ _1692_ _1694_ _1903_ net120 VGND VGND VPWR VPWR _1905_ sky130_fd_sc_hd__a211oi_4
X_5328_ _0756_ _0757_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5259_ _0446_ _0539_ _0682_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4630_ _3727_ _3728_ _3731_ _3587_ VGND VGND VPWR VPWR _3732_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4561_ _3642_ _3662_ _3663_ VGND VGND VPWR VPWR _3664_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6300_ _1818_ _1819_ VGND VGND VPWR VPWR _1820_ sky130_fd_sc_hd__xnor2_1
X_4492_ _3595_ VGND VGND VPWR VPWR _3596_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7280_ _2285_ _2890_ _0866_ VGND VGND VPWR VPWR _2891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6231_ _1641_ _1743_ _1744_ VGND VGND VPWR VPWR _1746_ sky130_fd_sc_hd__and3_2
XFILLER_0_100_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _1666_ _1667_ _1660_ VGND VGND VPWR VPWR _1670_ sky130_fd_sc_hd__a21o_1
X_5113_ _0392_ _0489_ _0522_ _0523_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__a211o_4
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _1431_ _1432_ VGND VGND VPWR VPWR _1595_ sky130_fd_sc_hd__and2b_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _0331_ _0400_ _0402_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__nor3_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6995_ _2579_ _2580_ VGND VGND VPWR VPWR _2581_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5946_ _1319_ _1433_ VGND VGND VPWR VPWR _1434_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5877_ _1355_ _1356_ _1184_ _1186_ VGND VGND VPWR VPWR _1358_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4828_ _0109_ _0111_ _0113_ _0211_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__o31a_1
XFILLER_0_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4759_ net178 _2642_ _2686_ _3242_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7478_ _3490_ _3591_ _3162_ _3104_ VGND VGND VPWR VPWR _3105_ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6429_ _1953_ _1960_ _0181_ VGND VGND VPWR VPWR _1961_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3992_ _0816_ _1133_ _1253_ _2850_ VGND VGND VPWR VPWR _2861_ sky130_fd_sc_hd__or4_1
X_6780_ _0172_ _0052_ _1745_ _1767_ VGND VGND VPWR VPWR _2345_ sky130_fd_sc_hd__and4_1
X_5800_ _1011_ _1014_ _1273_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5731_ _2149_ net36 net37 _2106_ VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5662_ _0975_ _1091_ _1121_ _1123_ VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__a211o_4
XFILLER_0_72_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4613_ _2980_ _3694_ _3696_ _3715_ VGND VGND VPWR VPWR _3716_ sky130_fd_sc_hd__a31o_1
X_5593_ _0906_ _0913_ VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7401_ _2836_ _2838_ VGND VGND VPWR VPWR _3025_ sky130_fd_sc_hd__and2b_1
XFILLER_0_143_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4544_ _3645_ _3531_ _2434_ _2106_ VGND VGND VPWR VPWR _3647_ sky130_fd_sc_hd__and4_1
X_7332_ _2943_ _2948_ VGND VGND VPWR VPWR _2949_ sky130_fd_sc_hd__xnor2_2
Xmax_cap110 net111 VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__buf_1
XFILLER_0_41_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap121 _1543_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__buf_1
XFILLER_0_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7263_ _0571_ _2062_ _2683_ VGND VGND VPWR VPWR _2874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4475_ _3575_ _3577_ VGND VGND VPWR VPWR _3579_ sky130_fd_sc_hd__nand2_1
X_6214_ _1725_ _1726_ _3430_ _2499_ VGND VGND VPWR VPWR _1727_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_40_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7194_ _2767_ _2798_ VGND VGND VPWR VPWR _2799_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6145_ _2313_ _2379_ _0720_ _0873_ VGND VGND VPWR VPWR _1651_ sky130_fd_sc_hd__and4_1
XFILLER_0_99_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6076_ _1573_ _1574_ _1554_ VGND VGND VPWR VPWR _1576_ sky130_fd_sc_hd__o21ai_2
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5027_ _3296_ _3298_ _3291_ _3292_ _0429_ _0199_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__mux4_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6978_ _2536_ _2537_ _2560_ _2561_ VGND VGND VPWR VPWR _2562_ sky130_fd_sc_hd__nand4_2
XFILLER_0_153_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5929_ _1394_ _1413_ _1414_ VGND VGND VPWR VPWR _1415_ sky130_fd_sc_hd__or3_4
XFILLER_0_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_591 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4260_ _3363_ _3364_ _3356_ VGND VGND VPWR VPWR _3366_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4191_ _3297_ _3129_ _0958_ VGND VGND VPWR VPWR _3298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6901_ _2446_ _2447_ _2476_ _2477_ VGND VGND VPWR VPWR _2479_ sky130_fd_sc_hd__a211o_1
XFILLER_0_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6832_ _2402_ VGND VGND VPWR VPWR _2403_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3975_ _2664_ VGND VGND VPWR VPWR _2675_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6763_ _2271_ _2268_ VGND VGND VPWR VPWR _2327_ sky130_fd_sc_hd__and2b_1
XFILLER_0_72_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5714_ _1074_ _1076_ _1178_ _1179_ VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6694_ _2250_ _2251_ VGND VGND VPWR VPWR _2252_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5645_ _0042_ _2773_ VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5576_ _1011_ _1027_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4527_ _2925_ _3533_ _3532_ _3530_ VGND VGND VPWR VPWR _3630_ sky130_fd_sc_hd__a22o_1
X_7315_ _2912_ _2929_ VGND VGND VPWR VPWR _2930_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4458_ _3558_ _3559_ _3560_ VGND VGND VPWR VPWR _3562_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_111_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7246_ _2854_ _2855_ VGND VGND VPWR VPWR _2856_ sky130_fd_sc_hd__xor2_1
X_7177_ _2578_ _2580_ VGND VGND VPWR VPWR _2780_ sky130_fd_sc_hd__or2_1
X_4389_ _3127_ _3493_ VGND VGND VPWR VPWR _3494_ sky130_fd_sc_hd__nand2_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6128_ _1384_ _1608_ _1483_ _1485_ VGND VGND VPWR VPWR _1632_ sky130_fd_sc_hd__a211oi_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _0281_ _1887_ VGND VGND VPWR VPWR _1557_ sky130_fd_sc_hd__and2_1
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3760_ _0314_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__buf_6
XFILLER_0_27_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5430_ _3284_ _3729_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5361_ _0791_ _0792_ _0784_ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5292_ _0461_ _0669_ _0667_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__o21a_1
X_4312_ _0652_ _3392_ _3393_ _3417_ VGND VGND VPWR VPWR _3418_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7100_ _2051_ net56 VGND VGND VPWR VPWR _2695_ sky130_fd_sc_hd__and2_1
X_4243_ _3342_ _3348_ VGND VGND VPWR VPWR _3349_ sky130_fd_sc_hd__xor2_4
XFILLER_0_10_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7031_ _2618_ _2619_ VGND VGND VPWR VPWR _2621_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4174_ _3202_ _3216_ _3199_ VGND VGND VPWR VPWR _3281_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6815_ _2609_ _2382_ _2383_ VGND VGND VPWR VPWR _2384_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_65_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6746_ _2263_ _1821_ VGND VGND VPWR VPWR _2308_ sky130_fd_sc_hd__and2b_1
X_3958_ net8 VGND VGND VPWR VPWR _2489_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3889_ _1712_ _1723_ VGND VGND VPWR VPWR _1734_ sky130_fd_sc_hd__nor2_2
XFILLER_0_18_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6677_ _2194_ _2195_ _2231_ _2232_ VGND VGND VPWR VPWR _2233_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_45_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5628_ _1071_ _1072_ _1085_ VGND VGND VPWR VPWR _1086_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5559_ _1876_ _1008_ VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7229_ _2824_ _2584_ _2835_ VGND VGND VPWR VPWR _2837_ sky130_fd_sc_hd__and3_1
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_754 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4930_ _1002_ _0293_ _0218_ _0217_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__a31o_1
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4861_ _2881_ _0247_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6600_ _2140_ _2141_ _2146_ VGND VGND VPWR VPWR _2148_ sky130_fd_sc_hd__a21o_1
X_3812_ _0881_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__buf_4
XFILLER_0_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4792_ _0100_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_16_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_16 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3743_ _0063_ _0117_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__nor2_1
X_6531_ _2270_ _0293_ _1890_ _2072_ VGND VGND VPWR VPWR _2074_ sky130_fd_sc_hd__a31o_1
XFILLER_0_125_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6462_ _1853_ _1855_ _1852_ VGND VGND VPWR VPWR _1998_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput101 net101 VGND VGND VPWR VPWR zero_flag sky130_fd_sc_hd__buf_8
X_5413_ _3589_ _0826_ _0000_ VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_3_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6393_ _1922_ _1921_ VGND VGND VPWR VPWR _1923_ sky130_fd_sc_hd__or2_4
XFILLER_0_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5344_ _0774_ _0775_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__nor2_2
XFILLER_0_88_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5275_ _3132_ _3151_ _1100_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__mux2_1
X_4226_ _3331_ _3332_ VGND VGND VPWR VPWR _3333_ sky130_fd_sc_hd__and2b_1
X_7014_ _2599_ _2600_ _2586_ VGND VGND VPWR VPWR _2602_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_10_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4157_ _0630_ _0641_ VGND VGND VPWR VPWR _3265_ sky130_fd_sc_hd__or2_2
X_4088_ _3195_ VGND VGND VPWR VPWR _3196_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_148_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6729_ _1277_ _2289_ _2278_ VGND VGND VPWR VPWR _2290_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_151_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput14 A[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_2
Xinput25 A[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_4
XFILLER_0_154_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput36 B[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput47 B[22] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_4
Xinput58 B[3] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_6
XFILLER_0_149_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5060_ _0351_ _0350_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__or2b_1
X_4011_ _2346_ _1034_ _1023_ _1045_ _0958_ _0925_ VGND VGND VPWR VPWR _3066_ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5962_ _1963_ _1448_ VGND VGND VPWR VPWR _1451_ sky130_fd_sc_hd__nand2_2
X_4913_ _3213_ _0305_ _3301_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5893_ _2215_ _3620_ _1204_ _1203_ VGND VGND VPWR VPWR _1376_ sky130_fd_sc_hd__a31o_1
XFILLER_0_48_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4844_ _0228_ _0229_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4775_ _0119_ _0120_ _0153_ _0154_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__nor4_1
XFILLER_0_56_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6514_ _2052_ _2053_ _1990_ _1907_ VGND VGND VPWR VPWR _2055_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7494_ net82 net83 _3120_ _3121_ VGND VGND VPWR VPWR _3122_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6445_ _1969_ _1978_ VGND VGND VPWR VPWR _1979_ sky130_fd_sc_hd__xor2_1
X_6376_ _1886_ _1888_ _1902_ VGND VGND VPWR VPWR _1904_ sky130_fd_sc_hd__nor3_1
XFILLER_0_30_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5327_ _3644_ _2149_ _0104_ _0105_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__and4_1
XFILLER_0_11_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5258_ _0447_ _0408_ _0536_ _0537_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__a211oi_2
X_4209_ net55 net28 VGND VGND VPWR VPWR _3316_ sky130_fd_sc_hd__and2_1
X_5189_ _0604_ _0605_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_748 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_670 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4560_ _3659_ _3660_ _3661_ VGND VGND VPWR VPWR _3663_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4491_ _0783_ _0641_ VGND VGND VPWR VPWR _3595_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6230_ _1741_ _1742_ _1642_ _1584_ VGND VGND VPWR VPWR _1744_ sky130_fd_sc_hd__a211o_1
XFILLER_0_100_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ _1660_ _1666_ _1667_ VGND VGND VPWR VPWR _1669_ sky130_fd_sc_hd__nand3_1
X_5112_ _0519_ _0520_ _0501_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__a21oi_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6092_ _1473_ _1593_ VGND VGND VPWR VPWR _1594_ sky130_fd_sc_hd__xnor2_4
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _0403_ _0404_ _0405_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__nand3_2
XFILLER_0_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6994_ _2577_ _2578_ _2171_ _1008_ VGND VGND VPWR VPWR _2580_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_149_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5945_ _1431_ _1432_ VGND VGND VPWR VPWR _1433_ sky130_fd_sc_hd__xnor2_4
X_5876_ _1184_ _1186_ _1355_ _1356_ VGND VGND VPWR VPWR _1357_ sky130_fd_sc_hd__a211oi_2
X_4827_ _0103_ _0114_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4758_ _0281_ _3651_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4689_ _0057_ _0058_ _0059_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7477_ _2980_ _3100_ _3101_ _3103_ VGND VGND VPWR VPWR _3104_ sky130_fd_sc_hd__a31o_1
XFILLER_0_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6428_ _1930_ _1936_ _1959_ VGND VGND VPWR VPWR _1960_ sky130_fd_sc_hd__a21o_1
X_6359_ _1882_ _1883_ _1720_ _1851_ VGND VGND VPWR VPWR _1885_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_11_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3991_ _1657_ _1668_ _1679_ _1701_ _2839_ VGND VGND VPWR VPWR _2850_ sky130_fd_sc_hd__a32o_1
XFILLER_0_76_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5730_ _2106_ _2149_ _0339_ _0340_ VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__nand4_4
XFILLER_0_9_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5661_ _1119_ _1120_ _1101_ VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7400_ _2930_ _3022_ VGND VGND VPWR VPWR _3023_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4612_ _3701_ _3706_ _3708_ _3714_ VGND VGND VPWR VPWR _3715_ sky130_fd_sc_hd__or4_1
X_5592_ _1044_ _1046_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4543_ _0041_ _2434_ _3644_ _3645_ VGND VGND VPWR VPWR _3646_ sky130_fd_sc_hd__a22oi_2
X_7331_ _2944_ _2945_ _2946_ VGND VGND VPWR VPWR _2948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap122 _3370_ VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_102_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7262_ _2694_ _2872_ VGND VGND VPWR VPWR _2873_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6213_ _3271_ _2521_ _2565_ _3632_ VGND VGND VPWR VPWR _1726_ sky130_fd_sc_hd__a22oi_2
X_4474_ _3575_ _3577_ VGND VGND VPWR VPWR _3578_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7193_ _2768_ _2797_ VGND VGND VPWR VPWR _2798_ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6144_ _1648_ _1649_ VGND VGND VPWR VPWR _1650_ sky130_fd_sc_hd__xnor2_2
X_6075_ _1554_ _1573_ _1574_ VGND VGND VPWR VPWR _1575_ sky130_fd_sc_hd__or3_4
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5026_ _3087_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__clkbuf_4
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6977_ _2558_ _2559_ _2540_ VGND VGND VPWR VPWR _2561_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5928_ _1410_ _1411_ _1412_ VGND VGND VPWR VPWR _1414_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_48_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_700 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5859_ _1328_ _1337_ VGND VGND VPWR VPWR _1338_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_559 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_476 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4190_ _3135_ _2510_ _0903_ VGND VGND VPWR VPWR _3297_ sky130_fd_sc_hd__mux2_1
X_6900_ _2473_ _2474_ _2231_ _2233_ VGND VGND VPWR VPWR _2477_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6831_ _2390_ _2456_ _1169_ _1294_ VGND VGND VPWR VPWR _2402_ sky130_fd_sc_hd__and4_1
XFILLER_0_106_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3974_ _2653_ VGND VGND VPWR VPWR _2664_ sky130_fd_sc_hd__buf_4
XFILLER_0_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6762_ _2128_ _2273_ VGND VGND VPWR VPWR _2326_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5713_ _0095_ _0654_ _1175_ _1177_ VGND VGND VPWR VPWR _1179_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_17_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6693_ _2249_ net51 _1056_ _2246_ VGND VGND VPWR VPWR _2251_ sky130_fd_sc_hd__and4b_1
XFILLER_0_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5644_ _2532_ _1102_ _1103_ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_73_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5575_ _1011_ _1027_ VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7314_ _2916_ _2928_ VGND VGND VPWR VPWR _2929_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_142_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4526_ _0106_ _0215_ _3197_ _3272_ _3526_ VGND VGND VPWR VPWR _3629_ sky130_fd_sc_hd__a41o_2
XFILLER_0_41_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4457_ _3558_ _3559_ _3560_ VGND VGND VPWR VPWR _3561_ sky130_fd_sc_hd__or3_4
X_7245_ _2647_ _2649_ VGND VGND VPWR VPWR _2855_ sky130_fd_sc_hd__or2b_1
X_7176_ _2777_ _2778_ VGND VGND VPWR VPWR _2779_ sky130_fd_sc_hd__xor2_1
X_4388_ _3490_ _3145_ _3492_ _3108_ VGND VGND VPWR VPWR _3493_ sky130_fd_sc_hd__a211o_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6127_ _1483_ _1485_ _1384_ _1608_ VGND VGND VPWR VPWR _1631_ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ net178 net15 net16 _3242_ VGND VGND VPWR VPWR _1556_ sky130_fd_sc_hd__a22o_1
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5009_ net180 _0409_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__nand2_2
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5360_ _0784_ _0791_ _0792_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__nand3_2
XFILLER_0_2_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5291_ _0673_ _0675_ _0676_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__nor3b_1
X_4311_ _3398_ _3399_ _3416_ VGND VGND VPWR VPWR _3417_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4242_ _3346_ _3347_ VGND VGND VPWR VPWR _3348_ sky130_fd_sc_hd__or2_4
XFILLER_0_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7030_ _2617_ net54 _1002_ _2615_ VGND VGND VPWR VPWR _2619_ sky130_fd_sc_hd__and4b_1
X_4173_ _3276_ _3278_ _0652_ VGND VGND VPWR VPWR _3280_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6814_ _3513_ _2576_ _2609_ _3424_ VGND VGND VPWR VPWR _2383_ sky130_fd_sc_hd__a22o_1
X_3957_ _2357_ _2467_ _0936_ VGND VGND VPWR VPWR _2478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6745_ _2303_ _2306_ VGND VGND VPWR VPWR _2307_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3888_ _0587_ VGND VGND VPWR VPWR _1723_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6676_ _2229_ _2230_ _2196_ _2197_ VGND VGND VPWR VPWR _2232_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_33_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5627_ _1077_ _1084_ VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5558_ _1876_ _1008_ VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__nor2_1
X_4509_ _3559_ _3470_ _3611_ VGND VGND VPWR VPWR _3612_ sky130_fd_sc_hd__and3b_1
XFILLER_0_130_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5489_ net32 net64 _3537_ _3572_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__and4_1
X_7228_ _2824_ _2584_ _2835_ VGND VGND VPWR VPWR _2836_ sky130_fd_sc_hd__a21oi_2
X_7159_ _2553_ _2556_ _2758_ _2759_ VGND VGND VPWR VPWR _2760_ sky130_fd_sc_hd__a211o_1
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer70 _0680_ VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__buf_2
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4860_ net32 VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3811_ _0499_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4791_ _0079_ _0086_ _0170_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__or3_1
XANTENNA_17 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6530_ _2707_ _0100_ _3722_ VGND VGND VPWR VPWR _2072_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3742_ _0063_ _0117_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6461_ _1992_ _1993_ _1994_ VGND VGND VPWR VPWR _1997_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5412_ _0848_ _0850_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6392_ _1918_ _1919_ _1639_ VGND VGND VPWR VPWR _1922_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5343_ _3385_ _2215_ _0771_ _0773_ VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5274_ _0579_ _0570_ _0693_ _3596_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4225_ _3329_ _3330_ _3253_ _3255_ VGND VGND VPWR VPWR _3332_ sky130_fd_sc_hd__a211o_1
X_7013_ _2586_ _2599_ _2600_ VGND VGND VPWR VPWR _2601_ sky130_fd_sc_hd__and3_1
X_4156_ _2936_ _2958_ _3263_ VGND VGND VPWR VPWR _3264_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4087_ net61 VGND VGND VPWR VPWR _3195_ sky130_fd_sc_hd__buf_4
XFILLER_0_93_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4989_ _0377_ _0386_ _0387_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__nand3_1
XFILLER_0_108_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6728_ _0438_ _2279_ VGND VGND VPWR VPWR _2289_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6659_ _2211_ _2212_ VGND VGND VPWR VPWR _2213_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput37 B[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_2
Xinput15 A[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_4
Xinput26 A[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput48 B[23] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_4
Xinput59 B[4] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_6
XFILLER_0_52_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4010_ _3046_ _1428_ _0696_ VGND VGND VPWR VPWR _3056_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5961_ _1963_ _1448_ VGND VGND VPWR VPWR _1450_ sky130_fd_sc_hd__or2_2
XFILLER_0_149_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4912_ _3602_ _0304_ _3087_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5892_ _1372_ _1374_ VGND VGND VPWR VPWR _1375_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4843_ _0108_ _0109_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4774_ _0151_ _0152_ _0060_ _0121_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6513_ _1990_ _1907_ net200 _2053_ VGND VGND VPWR VPWR _2054_ sky130_fd_sc_hd__a211oi_4
X_7493_ net85 _3069_ _3074_ _3081_ VGND VGND VPWR VPWR _3121_ sky130_fd_sc_hd__and4b_1
XFILLER_0_55_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6444_ _1800_ _1977_ VGND VGND VPWR VPWR _1978_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6375_ _1886_ _1888_ _1902_ VGND VGND VPWR VPWR _1903_ sky130_fd_sc_hd__o21a_2
XFILLER_0_11_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5326_ _0247_ _0104_ _3512_ _3644_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_11_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5257_ _0679_ _0680_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__or2b_1
XFILLER_0_139_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4208_ _3311_ _3314_ VGND VGND VPWR VPWR _3315_ sky130_fd_sc_hd__xnor2_2
X_5188_ _0475_ _0476_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__and2_1
X_4139_ _3175_ _3178_ _3177_ VGND VGND VPWR VPWR _3247_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_98_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4490_ _3194_ _3573_ _3574_ _3414_ _3593_ VGND VGND VPWR VPWR _3594_ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6160_ _1664_ _1665_ _1661_ VGND VGND VPWR VPWR _1667_ sky130_fd_sc_hd__a21o_1
X_5111_ _0501_ _0519_ _0520_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__and3_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _1590_ _1591_ VGND VGND VPWR VPWR _1593_ sky130_fd_sc_hd__xor2_4
XFILLER_0_0_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _0411_ _0408_ _0409_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__and3b_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6993_ _2171_ _1008_ _2577_ _2578_ VGND VGND VPWR VPWR _2579_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_149_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5944_ _1157_ _1259_ _1258_ VGND VGND VPWR VPWR _1432_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_47_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5875_ _1353_ _1354_ _1213_ _1215_ VGND VGND VPWR VPWR _1356_ sky130_fd_sc_hd__a211oi_2
X_4826_ _0208_ _0209_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4757_ _0131_ _0134_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__xnor2_2
X_4688_ _0057_ _0058_ _0059_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__nand3_4
X_7476_ _0379_ _0543_ _3102_ VGND VGND VPWR VPWR _3103_ sky130_fd_sc_hd__o21a_1
XFILLER_0_70_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6427_ _1797_ _1778_ VGND VGND VPWR VPWR _1959_ sky130_fd_sc_hd__and2b_1
XFILLER_0_101_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6358_ _1720_ _1851_ _1882_ _1883_ VGND VGND VPWR VPWR _1884_ sky130_fd_sc_hd__o211a_4
X_5309_ _0723_ _0736_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6289_ _1806_ _1807_ VGND VGND VPWR VPWR _1808_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3990_ _0063_ net25 _0783_ _1734_ _2828_ VGND VGND VPWR VPWR _2839_ sky130_fd_sc_hd__a41o_1
XFILLER_0_128_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5660_ _1101_ _1119_ _1120_ VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__nor3_4
XFILLER_0_73_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4611_ _3194_ _3709_ _3710_ _3686_ _3713_ VGND VGND VPWR VPWR _3714_ sky130_fd_sc_hd__a221o_1
XFILLER_0_154_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5591_ _0904_ _1043_ VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__and2_1
XFILLER_0_142_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4542_ _3169_ VGND VGND VPWR VPWR _3645_ sky130_fd_sc_hd__buf_4
X_7330_ _2730_ _2731_ _2732_ VGND VGND VPWR VPWR _2946_ sky130_fd_sc_hd__or3_1
XFILLER_0_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap112 _0803_ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__buf_1
Xmax_cap123 _1176_ VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_2
X_4473_ _3482_ _3497_ _3576_ VGND VGND VPWR VPWR _3577_ sky130_fd_sc_hd__a21o_1
X_7261_ _0438_ _2871_ _1277_ VGND VGND VPWR VPWR _2872_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6212_ _3195_ _3431_ net9 net10 VGND VGND VPWR VPWR _1725_ sky130_fd_sc_hd__and4_1
XFILLER_0_40_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7192_ _2785_ _2796_ VGND VGND VPWR VPWR _2797_ sky130_fd_sc_hd__xnor2_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6143_ _1056_ net48 VGND VGND VPWR VPWR _1649_ sky130_fd_sc_hd__nand2_1
X_6074_ _1569_ _1571_ _1572_ VGND VGND VPWR VPWR _1574_ sky130_fd_sc_hd__a21oi_2
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5025_ _3727_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__buf_2
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6976_ _2540_ _2558_ _2559_ VGND VGND VPWR VPWR _2560_ sky130_fd_sc_hd__or3_2
XFILLER_0_67_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5927_ _1410_ _1411_ _1412_ VGND VGND VPWR VPWR _1413_ sky130_fd_sc_hd__and3_2
XFILLER_0_119_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5858_ _1335_ _1336_ VGND VGND VPWR VPWR _1337_ sky130_fd_sc_hd__xor2_4
XFILLER_0_134_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4809_ _0176_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5789_ _1260_ _1261_ VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__nor2_4
XFILLER_0_17_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7459_ _3127_ net25 _0783_ _1734_ _3084_ VGND VGND VPWR VPWR _3085_ sky130_fd_sc_hd__a41o_1
XFILLER_0_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_801 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_552 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6830_ _2456_ _1170_ _1295_ _2390_ VGND VGND VPWR VPWR _2400_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6761_ _3571_ _2310_ _2311_ _2323_ VGND VGND VPWR VPWR _2325_ sky130_fd_sc_hd__a31o_1
XFILLER_0_147_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3973_ _2642_ VGND VGND VPWR VPWR _2653_ sky130_fd_sc_hd__buf_6
X_5712_ _1175_ _1177_ _0095_ _0654_ VGND VGND VPWR VPWR _1178_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_9_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6692_ _1056_ net51 _2247_ _2249_ VGND VGND VPWR VPWR _2250_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_45_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5643_ _0373_ net8 net9 _3352_ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5574_ _0826_ _0836_ _0877_ _0887_ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_142_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4525_ _3529_ _3548_ _3549_ VGND VGND VPWR VPWR _3628_ sky130_fd_sc_hd__nand3_1
XFILLER_0_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7313_ _2919_ _2927_ VGND VGND VPWR VPWR _2928_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4456_ _3377_ _3471_ _3470_ VGND VGND VPWR VPWR _3560_ sky130_fd_sc_hd__a21o_1
X_7244_ _2852_ _2853_ VGND VGND VPWR VPWR _2854_ sky130_fd_sc_hd__and2b_1
X_4387_ _0980_ _3148_ VGND VGND VPWR VPWR _3492_ sky130_fd_sc_hd__nor2_1
X_7175_ _2226_ _1008_ VGND VGND VPWR VPWR _2778_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6126_ _1488_ _1497_ VGND VGND VPWR VPWR _1630_ sky130_fd_sc_hd__or2_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6057_ _0488_ _0390_ net15 net16 VGND VGND VPWR VPWR _1555_ sky130_fd_sc_hd__nand4_1
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5008_ _0406_ _0407_ _0208_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__o21ai_1
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6959_ _2355_ _2363_ _2362_ VGND VGND VPWR VPWR _2541_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5290_ _0686_ _0687_ _0698_ _0716_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__o211ai_4
X_4310_ _3406_ _3411_ _3413_ _3415_ VGND VGND VPWR VPWR _3416_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4241_ _3344_ _3345_ net1 net63 VGND VGND VPWR VPWR _3347_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_77_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4172_ _3276_ _3278_ VGND VGND VPWR VPWR _3279_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6813_ _3424_ _3512_ _2576_ VGND VGND VPWR VPWR _2382_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3956_ _2412_ _2456_ _2029_ VGND VGND VPWR VPWR _2467_ sky130_fd_sc_hd__mux2_4
XFILLER_0_58_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6744_ _1614_ _1955_ _2304_ _2305_ _2278_ VGND VGND VPWR VPWR _2306_ sky130_fd_sc_hd__a32o_1
XFILLER_0_147_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6675_ _2196_ _2197_ _2229_ _2230_ VGND VGND VPWR VPWR _2231_ sky130_fd_sc_hd__a211o_2
XFILLER_0_18_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3887_ _0554_ VGND VGND VPWR VPWR _1712_ sky130_fd_sc_hd__clkbuf_4
X_5626_ _1082_ _1083_ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__xor2_1
XFILLER_0_60_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5557_ _1007_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4508_ _3508_ net144 _3557_ VGND VGND VPWR VPWR _3611_ sky130_fd_sc_hd__nand3_2
XFILLER_0_112_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5488_ _0104_ _3537_ _0105_ _2149_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__a22oi_1
X_4439_ _3540_ _3541_ _3542_ VGND VGND VPWR VPWR _3543_ sky130_fd_sc_hd__nand3_2
X_7227_ _2825_ _2834_ VGND VGND VPWR VPWR _2835_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7158_ _2742_ _2743_ _2757_ VGND VGND VPWR VPWR _2759_ sky130_fd_sc_hd__nor3_2
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7089_ _2683_ _3161_ VGND VGND VPWR VPWR _2684_ sky130_fd_sc_hd__and2b_1
X_6109_ _1609_ _1610_ VGND VGND VPWR VPWR _1611_ sky130_fd_sc_hd__nor2_1
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer60 _3371_ VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_1
Xrebuffer71 _3178_ VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4790_ _0079_ _0086_ _0170_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3810_ _0183_ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__buf_2
XFILLER_0_68_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3741_ _0106_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__buf_6
XFILLER_0_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_18 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6460_ _1992_ _1993_ _1994_ VGND VGND VPWR VPWR _1995_ sky130_fd_sc_hd__nand3_1
XFILLER_0_82_383 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5411_ _3212_ _3729_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__nand2_2
XFILLER_0_30_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6391_ _1639_ _1918_ _1919_ VGND VGND VPWR VPWR _1921_ sky130_fd_sc_hd__and3_1
X_5342_ _0771_ _0773_ _3631_ _2215_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_51_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7012_ _2427_ _2588_ _2597_ VGND VGND VPWR VPWR _2600_ sky130_fd_sc_hd__nand3_2
X_5273_ _0579_ _0570_ _0693_ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4224_ _3253_ _3255_ _3329_ _3330_ VGND VGND VPWR VPWR _3331_ sky130_fd_sc_hd__o211a_1
X_4155_ _2903_ _2335_ VGND VGND VPWR VPWR _3263_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4086_ net123 VGND VGND VPWR VPWR _3194_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4988_ _0383_ _0384_ _0385_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3939_ _2237_ _2270_ _2029_ VGND VGND VPWR VPWR _2281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6727_ _0861_ _3705_ _2287_ _3118_ VGND VGND VPWR VPWR _2288_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_614 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6658_ _2202_ _2210_ VGND VGND VPWR VPWR _2212_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5609_ _1037_ _1063_ _1064_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__nor3_2
XFILLER_0_143_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6589_ _2133_ _2134_ _2135_ VGND VGND VPWR VPWR _2136_ sky130_fd_sc_hd__nand3_1
XFILLER_0_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput27 A[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_8
Xinput16 A[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_4
XFILLER_0_107_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_832 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput49 B[24] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_2
Xinput38 B[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_4
XFILLER_0_52_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5960_ net48 VGND VGND VPWR VPWR _1448_ sky130_fd_sc_hd__clkbuf_4
X_5891_ _1370_ _1371_ _3709_ VGND VGND VPWR VPWR _1374_ sky130_fd_sc_hd__a21oi_1
X_4911_ _3134_ _3133_ _2675_ _3137_ _3046_ _3591_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__mux4_2
XFILLER_0_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_717 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4842_ _0225_ _0227_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4773_ _0060_ _0121_ _0151_ _0152_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_117_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_692 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6512_ _2025_ _2026_ _2049_ _2050_ VGND VGND VPWR VPWR _2053_ sky130_fd_sc_hd__o22a_1
X_7492_ net78 net79 net81 _3119_ VGND VGND VPWR VPWR _3120_ sky130_fd_sc_hd__nor4_2
XFILLER_0_55_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6443_ _1970_ _1976_ VGND VGND VPWR VPWR _1977_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_141_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6374_ _1893_ _1901_ VGND VGND VPWR VPWR _1902_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5325_ _3530_ _0110_ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__nand2_1
X_5256_ _0677_ _0678_ _0533_ _0536_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__a211o_1
XFILLER_0_54_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4207_ _3312_ _3313_ VGND VGND VPWR VPWR _3314_ sky130_fd_sc_hd__and2b_1
X_5187_ _0602_ _0603_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__nor2_2
X_4138_ _3243_ _3244_ _3241_ VGND VGND VPWR VPWR _3246_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4069_ net194 net44 net28 net33 VGND VGND VPWR VPWR _3178_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_504 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5110_ _0516_ _0517_ _0518_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__a21o_1
X_6090_ _1323_ _1427_ _1426_ VGND VGND VPWR VPWR _1591_ sky130_fd_sc_hd__o21ba_2
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _0320_ _0418_ _0444_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__a21o_2
XFILLER_0_85_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6992_ _2226_ _2270_ _0721_ _0874_ VGND VGND VPWR VPWR _2578_ sky130_fd_sc_hd__and4_1
XFILLER_0_149_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5943_ _1429_ _1430_ VGND VGND VPWR VPWR _1431_ sky130_fd_sc_hd__nand2_4
XFILLER_0_75_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5874_ _1213_ _1215_ _1353_ _1354_ VGND VGND VPWR VPWR _1355_ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4825_ _0102_ _0116_ _0119_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__or3_1
XFILLER_0_16_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4756_ _0132_ _0133_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_640 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4687_ _3649_ _3658_ _3657_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__a21bo_1
X_7475_ _0379_ _0543_ _3265_ VGND VGND VPWR VPWR _3102_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6426_ _1954_ _1956_ _1953_ VGND VGND VPWR VPWR _1958_ sky130_fd_sc_hd__a21o_1
X_6357_ _1870_ _1871_ _1881_ VGND VGND VPWR VPWR _1883_ sky130_fd_sc_hd__o21ai_2
X_5308_ _0734_ _0735_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6288_ _1794_ _1795_ _1804_ VGND VGND VPWR VPWR _1807_ sky130_fd_sc_hd__a21oi_1
X_5239_ _0470_ _0653_ _0659_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__or3_1
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4610_ _3712_ _3686_ VGND VGND VPWR VPWR _3713_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5590_ _0904_ _1043_ VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__nor2_1
X_4541_ net31 VGND VGND VPWR VPWR _3644_ sky130_fd_sc_hd__buf_4
XFILLER_0_53_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap113 _0648_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_1
Xmax_cap124 _3158_ VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
X_4472_ _3425_ _2182_ VGND VGND VPWR VPWR _3576_ sky130_fd_sc_hd__and2b_1
XFILLER_0_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7260_ _2051_ net56 VGND VGND VPWR VPWR _2871_ sky130_fd_sc_hd__nand2_1
Xmax_cap102 _2849_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__buf_1
X_6211_ _2892_ _2576_ _1565_ _1564_ _1865_ VGND VGND VPWR VPWR _1724_ sky130_fd_sc_hd__a32o_2
X_7191_ _2793_ _2794_ VGND VGND VPWR VPWR _2796_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6142_ _1645_ _1647_ VGND VGND VPWR VPWR _1648_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _1569_ _1571_ _1572_ VGND VGND VPWR VPWR _1573_ sky130_fd_sc_hd__and3_2
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _0422_ _0426_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__xnor2_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6975_ _2556_ _2557_ _2541_ VGND VGND VPWR VPWR _2559_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5926_ _1232_ _1240_ _1239_ VGND VGND VPWR VPWR _1412_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5857_ _1160_ _1163_ VGND VGND VPWR VPWR _1336_ sky130_fd_sc_hd__or2_2
XFILLER_0_17_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4808_ _2707_ _0100_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__and2_1
X_5788_ _1258_ _1259_ _1157_ VGND VGND VPWR VPWR _1261_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4739_ _0103_ _0114_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_50_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7458_ _0885_ _3083_ _0838_ VGND VGND VPWR VPWR _3084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6409_ _0187_ _0710_ _1283_ _1939_ _0429_ _0189_ VGND VGND VPWR VPWR _1940_ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7389_ _3008_ _3010_ VGND VGND VPWR VPWR _3011_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xsplit54 _3176_ VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_82_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6760_ _0844_ _2315_ _2318_ _2322_ VGND VGND VPWR VPWR _2323_ sky130_fd_sc_hd__a211o_1
X_3972_ net4 VGND VGND VPWR VPWR _2642_ sky130_fd_sc_hd__buf_4
XFILLER_0_85_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5711_ _3442_ _0326_ _0453_ _3635_ VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_57_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6691_ _0215_ _0346_ _1607_ net50 VGND VGND VPWR VPWR _2249_ sky130_fd_sc_hd__and4_1
XFILLER_0_45_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5642_ _3352_ _0373_ net8 VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5573_ _2095_ _0578_ _1020_ _1025_ VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__a211o_1
XFILLER_0_14_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4524_ _3615_ _3626_ VGND VGND VPWR VPWR _3627_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7312_ _2922_ _2926_ VGND VGND VPWR VPWR _2927_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4455_ net144 _3557_ _3508_ VGND VGND VPWR VPWR _3559_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_111_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7243_ net197 _2851_ _2610_ _2651_ VGND VGND VPWR VPWR _2853_ sky130_fd_sc_hd__o211ai_1
X_4386_ _3132_ _3138_ _3151_ _3136_ _1723_ _3490_ VGND VGND VPWR VPWR _3491_ sky130_fd_sc_hd__mux4_1
X_7174_ _2775_ _2776_ VGND VGND VPWR VPWR _2777_ sky130_fd_sc_hd__nand2_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6125_ _1495_ _1496_ VGND VGND VPWR VPWR _1629_ sky130_fd_sc_hd__or2b_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _1544_ _1553_ VGND VGND VPWR VPWR _1554_ sky130_fd_sc_hd__xnor2_2
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5007_ _0208_ _0406_ _0407_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__or3_4
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6958_ _2381_ _2538_ _2539_ VGND VGND VPWR VPWR _2540_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5909_ _1391_ _1392_ VGND VGND VPWR VPWR _1393_ sky130_fd_sc_hd__and2b_1
XFILLER_0_64_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6889_ _2457_ _2464_ VGND VGND VPWR VPWR _2465_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4240_ net1 _3343_ _3344_ _3345_ VGND VGND VPWR VPWR _3346_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_77_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4171_ _3215_ _3264_ _3277_ VGND VGND VPWR VPWR _3278_ sky130_fd_sc_hd__a21o_1
XFILLER_0_93_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6812_ _2377_ _2380_ VGND VGND VPWR VPWR _2381_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3955_ _2445_ VGND VGND VPWR VPWR _2456_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6743_ _1950_ _1954_ _2279_ _2119_ VGND VGND VPWR VPWR _2305_ sky130_fd_sc_hd__o211ai_1
X_6674_ _2227_ _2228_ _2213_ VGND VGND VPWR VPWR _2230_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_46_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3886_ _1690_ VGND VGND VPWR VPWR _1701_ sky130_fd_sc_hd__buf_2
X_5625_ _0934_ _0935_ VGND VGND VPWR VPWR _1083_ sky130_fd_sc_hd__nor2_2
XFILLER_0_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5556_ net45 VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__clkbuf_4
X_4507_ _3479_ _3567_ _3566_ VGND VGND VPWR VPWR _3610_ sky130_fd_sc_hd__o21ba_4
X_5487_ _0930_ _0931_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4438_ _3447_ _3450_ _3453_ VGND VGND VPWR VPWR _3542_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_111_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7226_ _2826_ _2833_ VGND VGND VPWR VPWR _2834_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4369_ net146 _3334_ _3378_ _3473_ VGND VGND VPWR VPWR _3474_ sky130_fd_sc_hd__o31ai_1
X_7157_ _2742_ _2743_ _2757_ VGND VGND VPWR VPWR _2758_ sky130_fd_sc_hd__o21a_2
XFILLER_0_10_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7088_ _0848_ _0196_ VGND VGND VPWR VPWR _2683_ sky130_fd_sc_hd__nor2_1
X_6108_ _1756_ _1608_ VGND VGND VPWR VPWR _1610_ sky130_fd_sc_hd__and2_1
X_6039_ _1532_ _1533_ _1529_ _1372_ VGND VGND VPWR VPWR _1535_ sky130_fd_sc_hd__a211o_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer72 _3376_ VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer50 _1921_ VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_1
Xrebuffer61 _1915_ VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_383 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3740_ _0095_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__buf_6
XFILLER_0_7_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_19 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_395 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5410_ _0428_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__buf_2
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6390_ _1916_ _1917_ _1790_ _1746_ VGND VGND VPWR VPWR _1919_ sky130_fd_sc_hd__a211o_1
XFILLER_0_140_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5341_ _3632_ _3271_ _3651_ _0491_ VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7011_ _2427_ _2588_ _2597_ VGND VGND VPWR VPWR _2599_ sky130_fd_sc_hd__a21o_1
X_5272_ _3571_ _0697_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__nand2_2
X_4223_ _3327_ _3328_ _3310_ VGND VGND VPWR VPWR _3330_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4154_ _3191_ net176 _3260_ VGND VGND VPWR VPWR _3262_ sky130_fd_sc_hd__nand3_1
XFILLER_0_128_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4085_ _0652_ _2969_ _3167_ _3193_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__a211o_2
XFILLER_0_148_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4987_ _0383_ _0384_ _0385_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__nand3_1
XFILLER_0_74_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6726_ _0861_ _2286_ VGND VGND VPWR VPWR _2287_ sky130_fd_sc_hd__nor2_1
X_3938_ _2259_ VGND VGND VPWR VPWR _2270_ sky130_fd_sc_hd__buf_4
XFILLER_0_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3869_ _1417_ _1439_ _1504_ VGND VGND VPWR VPWR _1515_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6657_ _2202_ _2210_ VGND VGND VPWR VPWR _2211_ sky130_fd_sc_hd__or2_1
XFILLER_0_143_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6588_ _0303_ _1767_ VGND VGND VPWR VPWR _2135_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5608_ _1061_ _1062_ _0942_ _1038_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5539_ net106 _0987_ _0806_ _0808_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7209_ _2813_ _2814_ VGND VGND VPWR VPWR _2815_ sky130_fd_sc_hd__or2_1
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput28 A[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_4
XFILLER_0_91_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput17 A[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_4
XFILLER_0_80_844 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput39 B[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_2
XFILLER_0_40_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5890_ _3709_ _1370_ _1371_ VGND VGND VPWR VPWR _1372_ sky130_fd_sc_hd__and3_1
X_4910_ _0175_ _0186_ _0296_ _3596_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_142_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4841_ _0205_ _0110_ _0223_ _0224_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_87_476 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4772_ _0148_ _0149_ _0130_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_117_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7491_ net75 net76 net77 _3117_ VGND VGND VPWR VPWR _3119_ sky130_fd_sc_hd__or4_4
XFILLER_0_71_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6511_ _2025_ _2026_ _2049_ _2050_ VGND VGND VPWR VPWR _2052_ sky130_fd_sc_hd__nor4_2
XFILLER_0_55_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6442_ _1973_ _1975_ VGND VGND VPWR VPWR _1976_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6373_ _1899_ _1900_ VGND VGND VPWR VPWR _1901_ sky130_fd_sc_hd__xor2_1
XFILLER_0_70_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5324_ _0752_ _0753_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5255_ _0533_ _0536_ _0677_ _0678_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__o211a_1
X_4206_ net58 _0074_ net26 net59 VGND VGND VPWR VPWR _3313_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5186_ _2379_ _0110_ _0600_ _0601_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__o2bb2a_1
X_4137_ _3241_ _3243_ _3244_ VGND VGND VPWR VPWR _3245_ sky130_fd_sc_hd__nand3_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4068_ net194 net33 _3176_ net28 VGND VGND VPWR VPWR _3177_ sky130_fd_sc_hd__nand4_2
XFILLER_0_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6709_ _2240_ _2267_ VGND VGND VPWR VPWR _2268_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _0419_ _0424_ _0425_ _0443_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__a31o_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6991_ _2270_ _0722_ _0875_ _2226_ VGND VGND VPWR VPWR _2577_ sky130_fd_sc_hd__a22oi_1
X_5942_ _1426_ _1427_ _1323_ VGND VGND VPWR VPWR _1430_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_146_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5873_ _1350_ _1352_ _1338_ VGND VGND VPWR VPWR _1354_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4824_ _0116_ _0119_ _0102_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4755_ _0161_ _3531_ net32 _3537_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__and4_1
XFILLER_0_56_671 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4686_ _0055_ _0056_ _0047_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__a21o_1
X_7474_ _0379_ _0728_ VGND VGND VPWR VPWR _3101_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6425_ _1953_ _1954_ _1956_ VGND VGND VPWR VPWR _1957_ sky130_fd_sc_hd__nand3_1
X_6356_ _1870_ _1871_ _1881_ VGND VGND VPWR VPWR _1882_ sky130_fd_sc_hd__or3_4
XFILLER_0_3_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5307_ _0664_ _0660_ _0661_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6287_ _1805_ VGND VGND VPWR VPWR _1806_ sky130_fd_sc_hd__inv_2
X_5238_ _0470_ _0653_ _0659_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5169_ _0558_ _3135_ _3134_ _3133_ _0583_ _0584_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_638 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4540_ _2881_ _2379_ VGND VGND VPWR VPWR _3643_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap114 _0398_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__buf_1
X_4471_ _3573_ _3574_ VGND VGND VPWR VPWR _3575_ sky130_fd_sc_hd__or2_2
XFILLER_0_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap103 _1989_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__buf_1
XFILLER_0_111_746 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6210_ _1546_ _1549_ VGND VGND VPWR VPWR _1722_ sky130_fd_sc_hd__nand2_1
X_7190_ _2589_ _2595_ _2594_ VGND VGND VPWR VPWR _2794_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6141_ _0215_ _1169_ _1294_ _0346_ VGND VGND VPWR VPWR _1647_ sky130_fd_sc_hd__a22o_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _1400_ _1409_ _1408_ VGND VGND VPWR VPWR _1572_ sky130_fd_sc_hd__a21bo_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _3134_ _0337_ _0300_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__a21oi_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6974_ _2541_ _2556_ _2557_ VGND VGND VPWR VPWR _2558_ sky130_fd_sc_hd__and3_1
X_5925_ _1408_ _1409_ _1400_ VGND VGND VPWR VPWR _1411_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5856_ _1333_ _1334_ VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__or2_2
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_747 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4807_ _3097_ _0188_ _0189_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5787_ _1157_ _1258_ _1259_ VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4738_ _0112_ _0113_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_16_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4669_ _0033_ _0038_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__xnor2_2
X_7457_ _3298_ _3300_ _3299_ _3082_ _0587_ _1712_ VGND VGND VPWR VPWR _3083_ sky130_fd_sc_hd__mux4_1
XFILLER_0_142_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6408_ _1778_ _1756_ _1963_ _1942_ _0583_ _0584_ VGND VGND VPWR VPWR _1939_ sky130_fd_sc_hd__mux4_1
XFILLER_0_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7388_ _2727_ _2735_ _3009_ VGND VGND VPWR VPWR _3010_ sky130_fd_sc_hd__a21oi_1
X_6339_ _1931_ _1861_ _1862_ VGND VGND VPWR VPWR _1863_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_99_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3971_ _2554_ _2620_ _0936_ VGND VGND VPWR VPWR _2631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5710_ _3635_ _3442_ _0325_ _0452_ VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__and4_1
XFILLER_0_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6690_ _2246_ VGND VGND VPWR VPWR _2247_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5641_ _1092_ _1099_ VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5572_ _0855_ _1009_ _1010_ _0854_ _1024_ VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4523_ _3624_ _3625_ VGND VGND VPWR VPWR _3626_ sky130_fd_sc_hd__or2_1
X_7311_ _2923_ _2924_ VGND VGND VPWR VPWR _2926_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7242_ _2610_ _2651_ net197 _2851_ VGND VGND VPWR VPWR _2852_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_40_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4454_ _3508_ _3556_ _3557_ VGND VGND VPWR VPWR _3558_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4385_ _1100_ VGND VGND VPWR VPWR _3490_ sky130_fd_sc_hd__clkbuf_4
X_7173_ _2270_ _2664_ _0722_ _0875_ VGND VGND VPWR VPWR _2776_ sky130_fd_sc_hd__nand4_1
XFILLER_0_1_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6124_ _1473_ _1593_ _1627_ VGND VGND VPWR VPWR _1628_ sky130_fd_sc_hd__a21bo_2
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _1551_ _1552_ VGND VGND VPWR VPWR _1553_ sky130_fd_sc_hd__and2b_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _0403_ _0404_ net179 VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__a21oi_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6957_ _2386_ _2387_ VGND VGND VPWR VPWR _2539_ sky130_fd_sc_hd__and2b_1
XFILLER_0_91_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5908_ _1389_ _1390_ _1386_ VGND VGND VPWR VPWR _1392_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6888_ _2462_ _2463_ VGND VGND VPWR VPWR _2464_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5839_ _0419_ _1306_ _1311_ _0573_ _1315_ VGND VGND VPWR VPWR _1316_ sky130_fd_sc_hd__a221o_1
XFILLER_0_134_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4170_ _3198_ _2412_ VGND VGND VPWR VPWR _3277_ sky130_fd_sc_hd__and2b_1
XFILLER_0_93_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6811_ _2376_ _2378_ _0295_ VGND VGND VPWR VPWR _2380_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3954_ _2434_ VGND VGND VPWR VPWR _2445_ sky130_fd_sc_hd__buf_4
XFILLER_0_46_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6742_ _1953_ _2280_ VGND VGND VPWR VPWR _2304_ sky130_fd_sc_hd__nor2_1
X_3885_ net68 net67 net66 VGND VGND VPWR VPWR _1690_ sky130_fd_sc_hd__and3b_1
XFILLER_0_58_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6673_ _2213_ _2227_ _2228_ VGND VGND VPWR VPWR _2229_ sky130_fd_sc_hd__and3_2
XFILLER_0_46_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5624_ _1080_ _1081_ VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5555_ _1006_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_4
X_4506_ _3561_ _3562_ _3563_ VGND VGND VPWR VPWR _3609_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5486_ _2324_ _0219_ _0928_ _0929_ VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4437_ _3538_ _3539_ _3536_ VGND VGND VPWR VPWR _3541_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7225_ _2831_ _2832_ VGND VGND VPWR VPWR _2833_ sky130_fd_sc_hd__nand2_1
X_7156_ _2748_ _2756_ VGND VGND VPWR VPWR _2757_ sky130_fd_sc_hd__xor2_1
Xwire4 _2052_ VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__buf_2
XFILLER_0_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4368_ _3374_ _3375_ _3376_ VGND VGND VPWR VPWR _3473_ sky130_fd_sc_hd__nand3_1
XFILLER_0_67_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6107_ _1756_ _1608_ VGND VGND VPWR VPWR _1609_ sky130_fd_sc_hd__nor2_1
X_4299_ _3127_ _3404_ VGND VGND VPWR VPWR _3405_ sky130_fd_sc_hd__nand2_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7087_ _1277_ _2680_ _2681_ VGND VGND VPWR VPWR _2682_ sky130_fd_sc_hd__o21a_1
X_6038_ _1529_ _1372_ _1532_ _1533_ VGND VGND VPWR VPWR _1534_ sky130_fd_sc_hd__o211ai_4
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer73 _0415_ VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer62 net210 VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_1
Xrebuffer40 _0552_ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer51 _1921_ VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__buf_1
XFILLER_0_139_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_831 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_395 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_638 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5340_ _3271_ _2248_ _0491_ _3196_ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5271_ _0693_ _0695_ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__xor2_1
X_4222_ _3310_ _3327_ _3328_ VGND VGND VPWR VPWR _3329_ sky130_fd_sc_hd__nand3_2
X_7010_ _2589_ _2596_ VGND VGND VPWR VPWR _2597_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4153_ _3259_ _3260_ _3191_ VGND VGND VPWR VPWR _3261_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4084_ _1657_ _3190_ _3191_ _3192_ VGND VGND VPWR VPWR _3193_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_144_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_614 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4986_ _0254_ _0255_ _0256_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3937_ _2248_ VGND VGND VPWR VPWR _2259_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6725_ _0433_ _0865_ _1466_ _2285_ _0866_ _0867_ VGND VGND VPWR VPWR _2286_ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3868_ _1449_ _1493_ VGND VGND VPWR VPWR _1504_ sky130_fd_sc_hd__xor2_1
XFILLER_0_61_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6656_ _2208_ _2209_ VGND VGND VPWR VPWR _2210_ sky130_fd_sc_hd__xor2_1
XFILLER_0_143_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6587_ _0401_ _1799_ net20 _0499_ VGND VGND VPWR VPWR _2134_ sky130_fd_sc_hd__a22o_1
X_3799_ _0303_ _0739_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__nand2_2
X_5607_ _0942_ _1038_ _1061_ _1062_ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_33_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5538_ _0806_ _0808_ net106 _0987_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_103_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5469_ _0909_ _0910_ _0751_ _0752_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__o211ai_1
X_7208_ _2812_ _2811_ VGND VGND VPWR VPWR _2814_ sky130_fd_sc_hd__and2b_1
X_7139_ _2725_ _2726_ _2736_ VGND VGND VPWR VPWR _2738_ sky130_fd_sc_hd__o21ai_2
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput18 A[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput29 A[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_4
XFILLER_0_91_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4840_ _0223_ _0224_ _1275_ _3619_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_87_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4771_ _0130_ _0148_ _0149_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__and3_1
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6510_ _2047_ _2048_ _2027_ _2028_ VGND VGND VPWR VPWR _2050_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7490_ net72 net73 net74 _3116_ VGND VGND VPWR VPWR _3117_ sky130_fd_sc_hd__or4_1
XFILLER_0_82_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6441_ _0991_ net51 _1971_ _1972_ VGND VGND VPWR VPWR _1975_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_140_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6372_ _3424_ _3512_ _2751_ _2773_ _1689_ VGND VGND VPWR VPWR _1900_ sky130_fd_sc_hd__a41o_1
XFILLER_0_71_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5323_ _0106_ _0220_ _0749_ _0751_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5254_ _0673_ _0675_ _0676_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__o21bai_1
X_4205_ net58 net59 net27 net26 VGND VGND VPWR VPWR _3312_ sky130_fd_sc_hd__and4_1
X_5185_ _0600_ _0601_ _2379_ _3619_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4136_ net44 net28 net29 net33 VGND VGND VPWR VPWR _3244_ sky130_fd_sc_hd__a22o_1
X_4067_ net44 VGND VGND VPWR VPWR _3176_ sky130_fd_sc_hd__buf_8
XFILLER_0_78_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4969_ _0361_ _0364_ _0365_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__nand3_1
XFILLER_0_47_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6708_ _1982_ _2266_ VGND VGND VPWR VPWR _2267_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6639_ net189 net104 _2189_ _2190_ VGND VGND VPWR VPWR _2191_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6990_ _2573_ _2574_ VGND VGND VPWR VPWR _2575_ sky130_fd_sc_hd__or2_1
X_5941_ _1323_ _1426_ _1427_ VGND VGND VPWR VPWR _1429_ sky130_fd_sc_hd__or3_1
XFILLER_0_88_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5872_ _1338_ _1350_ _1352_ VGND VGND VPWR VPWR _1353_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4823_ net150 _0076_ _0163_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__or3_1
XFILLER_0_118_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4754_ _0041_ _2149_ _2204_ _3645_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_90_439 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7473_ _0379_ _0728_ VGND VGND VPWR VPWR _3100_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4685_ _0047_ _0055_ _0056_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__nand3_2
XFILLER_0_114_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6424_ _1614_ _1955_ VGND VGND VPWR VPWR _1956_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6355_ _1872_ _1880_ VGND VGND VPWR VPWR _1881_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5306_ _0724_ _0733_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__xor2_2
XFILLER_0_59_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6286_ _1794_ _1795_ _1804_ VGND VGND VPWR VPWR _1805_ sky130_fd_sc_hd__nand3_2
X_5237_ _0655_ _0658_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__xor2_1
XFILLER_0_75_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5168_ _3591_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__clkbuf_4
X_5099_ _3448_ _0380_ _2489_ _3449_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4119_ _2062_ _3226_ _0587_ VGND VGND VPWR VPWR _3227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_530 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap115 net202 VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_2
X_4470_ _2237_ _3513_ VGND VGND VPWR VPWR _3574_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_758 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6140_ _0215_ _0346_ _1169_ _1294_ VGND VGND VPWR VPWR _1645_ sky130_fd_sc_hd__nand4_1
XFILLER_0_0_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _1562_ _1563_ _1568_ VGND VGND VPWR VPWR _1571_ sky130_fd_sc_hd__a21o_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _0295_ _0301_ _0422_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__a21o_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6973_ _2553_ _2555_ _2547_ VGND VGND VPWR VPWR _2557_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5924_ _1400_ _1408_ _1409_ VGND VGND VPWR VPWR _1410_ sky130_fd_sc_hd__nand3_1
XFILLER_0_152_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5855_ _0346_ net45 _1331_ _1332_ VGND VGND VPWR VPWR _1334_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4806_ _3301_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5786_ _1256_ _1257_ _1128_ _1158_ VGND VGND VPWR VPWR _1259_ sky130_fd_sc_hd__a211o_1
XFILLER_0_16_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4737_ _0021_ _0022_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4668_ _0034_ _0037_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__xor2_2
X_7456_ _1034_ _2346_ _1023_ _2412_ _0947_ _0914_ VGND VGND VPWR VPWR _3082_ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6407_ _1930_ _1936_ VGND VGND VPWR VPWR _1938_ sky130_fd_sc_hd__or2_1
XFILLER_0_141_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7387_ _2728_ _2734_ VGND VGND VPWR VPWR _3009_ sky130_fd_sc_hd__and2_1
X_4599_ _3137_ _2237_ _2182_ _2138_ _3046_ _3591_ VGND VGND VPWR VPWR _3702_ sky130_fd_sc_hd__mux4_1
XFILLER_0_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6338_ _0373_ _1887_ net15 _3352_ VGND VGND VPWR VPWR _1862_ sky130_fd_sc_hd__a22o_1
X_6269_ _1626_ _1753_ VGND VGND VPWR VPWR _1786_ sky130_fd_sc_hd__or2b_1
XFILLER_0_99_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xsplit67 _0030_ VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_66_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3970_ _2587_ _2609_ _2029_ VGND VGND VPWR VPWR _2620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5640_ _1093_ _1098_ VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5571_ _1009_ _1022_ VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4522_ _3515_ _3623_ VGND VGND VPWR VPWR _3625_ sky130_fd_sc_hd__nor2_1
X_7310_ _0328_ _0558_ VGND VGND VPWR VPWR _2924_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4453_ _3554_ _3555_ _3466_ _3468_ VGND VGND VPWR VPWR _3557_ sky130_fd_sc_hd__o211ai_4
X_7241_ _2802_ _2803_ _2847_ _2848_ VGND VGND VPWR VPWR _2851_ sky130_fd_sc_hd__o22a_1
XFILLER_0_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4384_ _3194_ _3480_ _3481_ _3414_ _3488_ VGND VGND VPWR VPWR _3489_ sky130_fd_sc_hd__a221o_1
X_7172_ _2664_ _0722_ _0875_ _2270_ VGND VGND VPWR VPWR _2775_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6123_ _1590_ _1591_ VGND VGND VPWR VPWR _1627_ sky130_fd_sc_hd__or2_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _1549_ _1550_ _1545_ VGND VGND VPWR VPWR _1552_ sky130_fd_sc_hd__a21o_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _0403_ _0404_ _0405_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6956_ _2387_ _2386_ VGND VGND VPWR VPWR _2538_ sky130_fd_sc_hd__or2b_1
XFILLER_0_49_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5907_ _1386_ _1389_ _1390_ VGND VGND VPWR VPWR _1391_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6887_ _2460_ _2461_ _2199_ _2201_ VGND VGND VPWR VPWR _2463_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_118_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5838_ _0861_ _3126_ _3213_ _1313_ _1314_ VGND VGND VPWR VPWR _1315_ sky130_fd_sc_hd__a311o_1
XFILLER_0_134_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5769_ _1236_ _1237_ _1238_ VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__a21o_1
XFILLER_0_91_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7439_ _2697_ _3063_ _2887_ _2883_ VGND VGND VPWR VPWR _3064_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_98_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6810_ _2375_ VGND VGND VPWR VPWR _2378_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3953_ _2423_ VGND VGND VPWR VPWR _2434_ sky130_fd_sc_hd__buf_6
XFILLER_0_9_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6741_ _2300_ _2301_ VGND VGND VPWR VPWR _2303_ sky130_fd_sc_hd__or2b_1
XFILLER_0_42_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3884_ _1570_ _1646_ VGND VGND VPWR VPWR _1679_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_523 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6672_ _2214_ _2216_ _2225_ VGND VGND VPWR VPWR _2228_ sky130_fd_sc_hd__nand3_1
XFILLER_0_46_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5623_ _2160_ _0110_ VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5554_ _0872_ _0894_ _1005_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__or3_1
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4505_ _3569_ _3570_ _3608_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__a21o_2
X_5485_ _2313_ net38 _0928_ _0929_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__nand4_2
X_4436_ _3536_ _3538_ _3539_ VGND VGND VPWR VPWR _3540_ sky130_fd_sc_hd__nand3_1
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7224_ _2827_ _2829_ _2830_ VGND VGND VPWR VPWR _2832_ sky130_fd_sc_hd__or3_1
X_4367_ _3470_ _3471_ VGND VGND VPWR VPWR _3472_ sky130_fd_sc_hd__or2b_1
X_7155_ _2754_ _2755_ VGND VGND VPWR VPWR _2756_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6106_ _1607_ VGND VGND VPWR VPWR _1608_ sky130_fd_sc_hd__clkbuf_4
X_4298_ _1723_ _3403_ VGND VGND VPWR VPWR _3404_ sky130_fd_sc_hd__nand2_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7086_ _2018_ net54 VGND VGND VPWR VPWR _2681_ sky130_fd_sc_hd__or2_1
X_6037_ _3620_ _2653_ _1530_ _1531_ VGND VGND VPWR VPWR _1533_ sky130_fd_sc_hd__a22o_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_818 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer30 _1422_ VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__buf_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer52 _3259_ VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_1
Xrebuffer41 net95 VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__buf_2
XFILLER_0_96_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer63 _1086_ VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__buf_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer74 _3374_ VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6939_ _2511_ _2512_ _2517_ VGND VGND VPWR VPWR _2519_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_843 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5270_ _0563_ _0567_ _0694_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4221_ _3324_ _3325_ _3326_ VGND VGND VPWR VPWR _3328_ sky130_fd_sc_hd__a21o_1
X_4152_ _1548_ _3189_ net211 _3258_ VGND VGND VPWR VPWR _3260_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_128_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4083_ _0783_ _1144_ _1154_ _1165_ VGND VGND VPWR VPWR _3192_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_78_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4985_ _0381_ _0382_ _0378_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3936_ net3 VGND VGND VPWR VPWR _2248_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6724_ _1821_ _1810_ _1778_ _1756_ _0863_ _0864_ VGND VGND VPWR VPWR _2285_ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3867_ _0750_ _1482_ VGND VGND VPWR VPWR _1493_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6655_ _2401_ _1007_ _2064_ _2063_ VGND VGND VPWR VPWR _2209_ sky130_fd_sc_hd__a31o_1
XFILLER_0_116_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6586_ _0499_ _0401_ _1799_ net20 VGND VGND VPWR VPWR _2133_ sky130_fd_sc_hd__nand4_1
X_3798_ _0324_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__buf_6
X_5606_ _1059_ _1060_ _1047_ VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__o21a_1
XFILLER_0_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5537_ _0921_ _0922_ _0984_ _0985_ VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__o22a_1
XFILLER_0_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5468_ _0751_ _0752_ _0909_ _0910_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7207_ _2811_ _2812_ VGND VGND VPWR VPWR _2813_ sky130_fd_sc_hd__and2b_1
XFILLER_0_111_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4419_ _0085_ _3433_ _3431_ _1264_ VGND VGND VPWR VPWR _3523_ sky130_fd_sc_hd__a22o_1
X_5399_ _0834_ _0835_ _0829_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_10_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7138_ _2725_ _2726_ _2736_ VGND VGND VPWR VPWR _2737_ sky130_fd_sc_hd__or3_2
X_7069_ _2660_ _2661_ VGND VGND VPWR VPWR _2662_ sky130_fd_sc_hd__nor2_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput19 A[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_2
XFILLER_0_135_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_670 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4770_ _0145_ _0146_ _0147_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__a21o_1
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6440_ _1971_ _1972_ _0991_ net51 VGND VGND VPWR VPWR _1973_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_140_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6371_ _1896_ _1897_ VGND VGND VPWR VPWR _1899_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5322_ _0095_ net38 _0749_ _0751_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__nand4_2
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5253_ _0673_ _0675_ _0676_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__or3b_1
X_4204_ _0324_ net60 VGND VGND VPWR VPWR _3311_ sky130_fd_sc_hd__nand2_1
X_5184_ _2423_ net31 net64 _3572_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__and4_1
X_4135_ _3242_ net44 net28 net29 VGND VGND VPWR VPWR _3243_ sky130_fd_sc_hd__nand4_2
X_4066_ _0281_ net26 VGND VGND VPWR VPWR _3175_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4968_ _3530_ _3385_ _0362_ _0363_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4899_ _0287_ _0289_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__nor2_1
X_3919_ _2051_ net25 _0892_ VGND VGND VPWR VPWR _2062_ sky130_fd_sc_hd__mux2_2
XFILLER_0_80_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6707_ _2241_ _2265_ VGND VGND VPWR VPWR _2266_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6638_ _2165_ _2166_ _2187_ _2188_ VGND VGND VPWR VPWR _2190_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_117_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6569_ _0304_ _0845_ _1308_ _2114_ _0866_ _0867_ VGND VGND VPWR VPWR _2115_ sky130_fd_sc_hd__mux4_1
XFILLER_0_100_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5940_ _1424_ _1425_ _1254_ net198 VGND VGND VPWR VPWR _1427_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5871_ _1180_ _1339_ _1349_ VGND VGND VPWR VPWR _1352_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4822_ _3305_ _0171_ _0173_ _0184_ _0206_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__a311o_4
XFILLER_0_75_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4753_ _2881_ _3644_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7472_ _3581_ _3584_ _3098_ _3582_ _0063_ _3301_ VGND VGND VPWR VPWR _3099_ sky130_fd_sc_hd__mux4_1
XFILLER_0_50_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4684_ _0051_ _0053_ _0054_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_723 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6423_ _1770_ _1930_ VGND VGND VPWR VPWR _1955_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6354_ _1873_ _1879_ VGND VGND VPWR VPWR _1880_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5305_ _0731_ _0732_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__and2_1
X_6285_ _1802_ _1803_ VGND VGND VPWR VPWR _1804_ sky130_fd_sc_hd__nand2_1
X_5236_ _0326_ _0656_ _0657_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_52_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5167_ _3046_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__clkbuf_4
X_5098_ _0292_ _2740_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__and2_1
X_4118_ _3224_ _3225_ _1712_ VGND VGND VPWR VPWR _3226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4049_ net66 net65 net68 net67 VGND VGND VPWR VPWR _3158_ sky130_fd_sc_hd__nor4b_2
XFILLER_0_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap116 _0155_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__buf_1
XFILLER_0_111_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap105 _1814_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__buf_1
XFILLER_0_151_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _1562_ _1563_ _1568_ VGND VGND VPWR VPWR _1569_ sky130_fd_sc_hd__nand3_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _0295_ _0301_ _0422_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__nand3_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6972_ _2547_ _2553_ _2555_ VGND VGND VPWR VPWR _2556_ sky130_fd_sc_hd__nand3_4
X_5923_ _1404_ _1405_ _1407_ VGND VGND VPWR VPWR _1409_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5854_ _0335_ net45 _1331_ _1332_ VGND VGND VPWR VPWR _1333_ sky130_fd_sc_hd__and4_1
XFILLER_0_8_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4805_ _3500_ _0187_ _3087_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5785_ _1128_ net199 _1256_ _1257_ VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_8_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4736_ _0109_ _0111_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4667_ _3635_ _0035_ _0036_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__a21bo_1
X_7455_ _3069_ _3074_ _3081_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__nand3_4
XFILLER_0_16_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7386_ _3720_ _0862_ VGND VGND VPWR VPWR _3008_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6406_ _1930_ _1936_ VGND VGND VPWR VPWR _1937_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6337_ _3352_ _0373_ _1887_ VGND VGND VPWR VPWR _1861_ sky130_fd_sc_hd__and3_1
X_4598_ _3580_ _3697_ _3700_ _3587_ VGND VGND VPWR VPWR _3701_ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6268_ _1785_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_6
X_5219_ _0636_ _0637_ _0628_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__a21o_1
X_6199_ _3169_ net191 net13 VGND VGND VPWR VPWR _1710_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5570_ _0438_ _1021_ _0000_ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__a21oi_1
X_4521_ _3515_ _3623_ VGND VGND VPWR VPWR _3624_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4452_ _3466_ _3468_ _3554_ _3555_ VGND VGND VPWR VPWR _3556_ sky130_fd_sc_hd__a211o_1
XFILLER_0_13_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7240_ _2802_ _2803_ _2847_ _2848_ VGND VGND VPWR VPWR _2849_ sky130_fd_sc_hd__nor4_1
XFILLER_0_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4383_ _3486_ _3487_ _3201_ VGND VGND VPWR VPWR _3488_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7171_ _2771_ _2772_ VGND VGND VPWR VPWR _2774_ sky130_fd_sc_hd__xor2_1
X_6122_ _1594_ _1596_ VGND VGND VPWR VPWR _1626_ sky130_fd_sc_hd__or2_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6053_ _1545_ _1549_ _1550_ VGND VGND VPWR VPWR _1551_ sky130_fd_sc_hd__and3_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _0210_ _0276_ _0275_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__a21bo_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6955_ _2534_ _2535_ _2353_ _2503_ VGND VGND VPWR VPWR _2537_ sky130_fd_sc_hd__a211o_1
XFILLER_0_119_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5906_ _3430_ _2740_ _1387_ _1388_ VGND VGND VPWR VPWR _1390_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6886_ _2199_ _2201_ _2460_ _2461_ VGND VGND VPWR VPWR _2462_ sky130_fd_sc_hd__a211o_1
XFILLER_0_118_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5837_ _0854_ _1297_ _1298_ _0855_ _1280_ VGND VGND VPWR VPWR _1314_ sky130_fd_sc_hd__a221o_1
XFILLER_0_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5768_ _1236_ _1237_ _1238_ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__nand3_1
XFILLER_0_63_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4719_ _0065_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5699_ _0434_ net45 _1161_ _1162_ VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__and4_1
XFILLER_0_16_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7438_ _2672_ _2677_ _2701_ VGND VGND VPWR VPWR _3063_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7369_ _2981_ _2988_ VGND VGND VPWR VPWR _2989_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_502 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6740_ _2007_ _2299_ VGND VGND VPWR VPWR _2301_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3952_ net30 VGND VGND VPWR VPWR _2423_ sky130_fd_sc_hd__buf_8
XFILLER_0_73_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3883_ _0783_ _1144_ _1154_ _1165_ VGND VGND VPWR VPWR _1668_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_73_535 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6671_ _2214_ _2216_ _2225_ VGND VGND VPWR VPWR _2227_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5622_ _3573_ _1079_ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5553_ _0320_ _0998_ _0999_ _1004_ VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4504_ _3571_ _3578_ _3579_ _3607_ VGND VGND VPWR VPWR _3608_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5484_ _3442_ _2434_ _0339_ _0340_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__nand4_4
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4435_ _3451_ _3452_ _2149_ _2204_ VGND VGND VPWR VPWR _3539_ sky130_fd_sc_hd__nand4_2
X_7223_ _2827_ _2829_ _2830_ VGND VGND VPWR VPWR _2831_ sky130_fd_sc_hd__o21ai_1
X_4366_ _3468_ _3469_ net183 _3419_ VGND VGND VPWR VPWR _3471_ sky130_fd_sc_hd__a211o_1
X_7154_ _2549_ _2551_ VGND VGND VPWR VPWR _2755_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6105_ net49 VGND VGND VPWR VPWR _1607_ sky130_fd_sc_hd__buf_2
X_4297_ _2073_ _1843_ _1712_ VGND VGND VPWR VPWR _3403_ sky130_fd_sc_hd__mux2_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7085_ _3589_ _2670_ VGND VGND VPWR VPWR _2680_ sky130_fd_sc_hd__nor2_1
X_6036_ _0110_ _2653_ _1530_ _1531_ VGND VGND VPWR VPWR _1532_ sky130_fd_sc_hd__nand4_4
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer20 _3556_ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__buf_6
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer31 _3628_ VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer64 _3379_ VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer53 _2111_ VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_1
Xrebuffer42 net87 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_139_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer75 _3257_ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6938_ _2511_ _2512_ _2517_ VGND VGND VPWR VPWR _2518_ sky130_fd_sc_hd__nand3_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6869_ _2191_ _2235_ VGND VGND VPWR VPWR _2443_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4220_ _3324_ _3325_ _3326_ VGND VGND VPWR VPWR _3327_ sky130_fd_sc_hd__nand3_2
X_4151_ _1548_ _3189_ net211 _3258_ VGND VGND VPWR VPWR _3259_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_49_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4082_ _1657_ _3189_ VGND VGND VPWR VPWR _3191_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4984_ _0378_ _0381_ _0382_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__nand3_1
X_3935_ _2226_ VGND VGND VPWR VPWR _2237_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6723_ _2282_ _2283_ VGND VGND VPWR VPWR _2284_ sky130_fd_sc_hd__or2_1
X_6654_ _2206_ _2207_ VGND VGND VPWR VPWR _2208_ sky130_fd_sc_hd__xor2_1
XFILLER_0_132_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3866_ _1460_ _1471_ VGND VGND VPWR VPWR _1482_ sky130_fd_sc_hd__and2b_1
X_5605_ _1047_ _1059_ _1060_ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__nor3_1
XFILLER_0_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3797_ _0685_ _0696_ _0717_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_82_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6585_ _2011_ _2012_ _2022_ VGND VGND VPWR VPWR _2132_ sky130_fd_sc_hd__nor3_2
XFILLER_0_14_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5536_ _0921_ _0922_ _0984_ _0985_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__nor4_1
XFILLER_0_41_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5467_ _0907_ _0908_ _0739_ net41 VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_111_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4418_ _2379_ _3443_ _3445_ _3441_ VGND VGND VPWR VPWR _3522_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_2_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7206_ _2617_ _2619_ VGND VGND VPWR VPWR _2812_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5398_ _0439_ _0425_ _0563_ _0693_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__a211o_1
X_4349_ _3447_ _3450_ _3453_ VGND VGND VPWR VPWR _3454_ sky130_fd_sc_hd__nand3_1
X_7137_ _2727_ _2735_ VGND VGND VPWR VPWR _2736_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7068_ _2483_ _2485_ _2659_ VGND VGND VPWR VPWR _2661_ sky130_fd_sc_hd__and3_1
X_6019_ _1498_ _1511_ _1512_ VGND VGND VPWR VPWR _1513_ sky130_fd_sc_hd__nand3_2
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_811 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6370_ _3619_ _2751_ VGND VGND VPWR VPWR _1897_ sky130_fd_sc_hd__and2_1
XFILLER_0_140_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5321_ _3635_ _3442_ _0339_ _0340_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__nand4_4
XFILLER_0_51_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5252_ _0463_ _0449_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__and2b_1
XFILLER_0_48_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4203_ _3306_ _3309_ VGND VGND VPWR VPWR _3310_ sky130_fd_sc_hd__xnor2_2
X_5183_ _2106_ _3422_ _0105_ _2434_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_48_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4134_ net33 VGND VGND VPWR VPWR _3242_ sky130_fd_sc_hd__buf_12
X_4065_ _3172_ _3173_ VGND VGND VPWR VPWR _3174_ sky130_fd_sc_hd__xor2_2
XFILLER_0_148_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4967_ _2445_ _3385_ _0362_ _0363_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__nand4_2
XFILLER_0_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4898_ _0086_ _0170_ _0288_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__a21bo_1
X_3918_ net24 VGND VGND VPWR VPWR _2051_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6706_ _2262_ _2264_ VGND VGND VPWR VPWR _2265_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3849_ _1275_ _0499_ _0401_ _0739_ VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__a22o_1
X_6637_ _2165_ _2166_ _2187_ _2188_ VGND VGND VPWR VPWR _2189_ sky130_fd_sc_hd__or4_4
XFILLER_0_62_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6568_ _1810_ _1778_ _1756_ _1963_ _0863_ _0864_ VGND VGND VPWR VPWR _2114_ sky130_fd_sc_hd__mux4_1
XFILLER_0_132_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5519_ _0964_ _0965_ _0963_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6499_ _3512_ _2499_ _2532_ _3423_ VGND VGND VPWR VPWR _2038_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5870_ _1180_ _1339_ _1349_ VGND VGND VPWR VPWR _1350_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_146_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4821_ _2980_ _0185_ _0186_ _0204_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__a31o_1
XFILLER_0_34_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4752_ _0122_ _0129_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4683_ _0051_ _0053_ _0054_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__nand3_1
X_7471_ _2467_ _3071_ _2193_ _2357_ _3077_ _0969_ VGND VGND VPWR VPWR _3098_ sky130_fd_sc_hd__mux4_1
XFILLER_0_50_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6422_ _1610_ _1929_ _1928_ VGND VGND VPWR VPWR _1954_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_44_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6353_ _1877_ _1878_ VGND VGND VPWR VPWR _1879_ sky130_fd_sc_hd__or2_4
XFILLER_0_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5304_ _0729_ _0730_ _0725_ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__o21ai_1
X_6284_ _1796_ _1801_ VGND VGND VPWR VPWR _1803_ sky130_fd_sc_hd__or2_1
X_5235_ _0324_ _0325_ _0453_ net163 VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5166_ _3414_ _0560_ _0561_ _3194_ _0581_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__a221o_1
X_5097_ _0502_ _0505_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__xnor2_2
X_4117_ _1974_ _1788_ _0947_ VGND VGND VPWR VPWR _3225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4048_ _3127_ _3141_ _3155_ _3156_ VGND VGND VPWR VPWR _3157_ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_0_149_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5999_ _1489_ _1490_ _0215_ net45 VGND VGND VPWR VPWR _1491_ sky130_fd_sc_hd__and4b_1
XFILLER_0_148_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_666 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap117 _2186_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__buf_1
XFILLER_0_52_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _0420_ _0421_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__or2_2
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6971_ _2550_ _2551_ _2552_ VGND VGND VPWR VPWR _2555_ sky130_fd_sc_hd__a21o_1
X_5922_ _1404_ _1405_ _1407_ VGND VGND VPWR VPWR _1408_ sky130_fd_sc_hd__nand3_1
XFILLER_0_76_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5853_ _3440_ _0720_ _0873_ _1275_ VGND VGND VPWR VPWR _1332_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5784_ net107 _1192_ _1254_ net205 VGND VGND VPWR VPWR _1257_ sky130_fd_sc_hd__o22ai_4
X_4804_ _3133_ _2675_ _3137_ _2237_ _3046_ _3591_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__mux4_2
XFILLER_0_29_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4735_ _0335_ _0110_ _0107_ _0108_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_8_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4666_ _2368_ _3433_ _3431_ _2302_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__a22o_1
X_7454_ _0860_ _3210_ _0196_ _3079_ _3080_ VGND VGND VPWR VPWR _3081_ sky130_fd_sc_hd__o311a_1
XFILLER_0_141_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7385_ _2903_ _1810_ VGND VGND VPWR VPWR _3007_ sky130_fd_sc_hd__nand2_1
X_4597_ _3127_ _3699_ VGND VGND VPWR VPWR _3700_ sky130_fd_sc_hd__nand2_1
X_6405_ _1770_ _1782_ _1935_ VGND VGND VPWR VPWR _1936_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6336_ _1856_ _1857_ _1858_ VGND VGND VPWR VPWR _1860_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6267_ _1617_ _1757_ _1769_ _1784_ VGND VGND VPWR VPWR _1785_ sky130_fd_sc_hd__or4_4
X_5218_ _0628_ _0636_ _0637_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__nand3_2
X_6198_ _1705_ _1706_ _1707_ VGND VGND VPWR VPWR _1709_ sky130_fd_sc_hd__a21o_1
X_5149_ _0562_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4520_ _3618_ _3622_ VGND VGND VPWR VPWR _3623_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4451_ _3552_ _3553_ _3519_ VGND VGND VPWR VPWR _3555_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_103_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7170_ _2456_ _1448_ VGND VGND VPWR VPWR _2772_ sky130_fd_sc_hd__nand2_1
X_4382_ _1100_ _0925_ _0969_ VGND VGND VPWR VPWR _3487_ sky130_fd_sc_hd__and3_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6121_ net153 _1620_ _1623_ VGND VGND VPWR VPWR _1625_ sky130_fd_sc_hd__and3_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6052_ _3430_ _2773_ _1546_ _1547_ VGND VGND VPWR VPWR _1550_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _0400_ _0402_ _0331_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__o21ai_2
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6954_ _2353_ _2503_ _2534_ _2535_ VGND VGND VPWR VPWR _2536_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_119_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5905_ _3631_ _2751_ _1387_ _1388_ VGND VGND VPWR VPWR _1389_ sky130_fd_sc_hd__nand4_1
XFILLER_0_146_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6885_ _2458_ _2459_ _0357_ _1949_ VGND VGND VPWR VPWR _2461_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_91_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5836_ _1298_ _1312_ VGND VGND VPWR VPWR _1313_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5767_ _1107_ _1109_ _1108_ VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_91_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4718_ _3624_ _0028_ _0091_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_115_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5698_ _1275_ _0720_ _0873_ _0739_ VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4649_ _3629_ _3641_ _3639_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7437_ _2672_ _2697_ VGND VGND VPWR VPWR _3062_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7368_ _2982_ _2987_ VGND VGND VPWR VPWR _2988_ sky130_fd_sc_hd__xnor2_1
X_7299_ _2907_ _2911_ VGND VGND VPWR VPWR _2912_ sky130_fd_sc_hd__xnor2_1
X_6319_ _1838_ _1839_ _1840_ VGND VGND VPWR VPWR _1841_ sky130_fd_sc_hd__nand3_1
XFILLER_0_87_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_831 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3951_ _2401_ VGND VGND VPWR VPWR _2412_ sky130_fd_sc_hd__buf_4
XFILLER_0_128_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3882_ _1570_ _1646_ VGND VGND VPWR VPWR _1657_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6670_ _2217_ _2224_ VGND VGND VPWR VPWR _2225_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5621_ _3422_ _3651_ VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5552_ _0878_ _1001_ _1003_ VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__o21a_1
XFILLER_0_53_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4503_ _3588_ _3594_ _3606_ VGND VGND VPWR VPWR _3607_ sky130_fd_sc_hd__or3b_1
XFILLER_0_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5483_ _2434_ net36 _0340_ _3442_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4434_ _3448_ net32 _3537_ _3449_ VGND VGND VPWR VPWR _3538_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7222_ _0117_ _1949_ VGND VGND VPWR VPWR _2830_ sky130_fd_sc_hd__nand2_1
X_4365_ net183 _3419_ _3468_ _3469_ VGND VGND VPWR VPWR _3470_ sky130_fd_sc_hd__o211a_1
X_7153_ _2752_ _2753_ VGND VGND VPWR VPWR _2754_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7084_ _2311_ _2672_ _2677_ _0181_ VGND VGND VPWR VPWR _2679_ sky130_fd_sc_hd__a31oi_1
X_6104_ _3571_ _1453_ _1455_ _1606_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__a31o_1
X_4296_ _3400_ _3401_ _0870_ VGND VGND VPWR VPWR _3402_ sky130_fd_sc_hd__mux2_1
X_6035_ _0105_ _2696_ _2740_ _0104_ VGND VGND VPWR VPWR _1531_ sky130_fd_sc_hd__a22o_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer21 _3257_ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_1
Xrebuffer10 _1135_ VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_1
Xrebuffer32 _0271_ VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__buf_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer54 _1437_ VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer43 net85 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_4
Xrebuffer76 _3670_ VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_89_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer65 _2025_ VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6937_ _2515_ _2516_ VGND VGND VPWR VPWR _2517_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6868_ _2440_ _2441_ VGND VGND VPWR VPWR _2442_ sky130_fd_sc_hd__and2b_1
XFILLER_0_9_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5819_ net47 VGND VGND VPWR VPWR _1294_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6799_ _2353_ _2354_ _2365_ VGND VGND VPWR VPWR _2366_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4150_ net160 _3256_ _3186_ _3231_ VGND VGND VPWR VPWR _3258_ sky130_fd_sc_hd__o211ai_1
Xoutput90 net90 VGND VGND VPWR VPWR result[29] sky130_fd_sc_hd__clkbuf_4
X_4081_ _1548_ _3189_ VGND VGND VPWR VPWR _3190_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4983_ _3451_ _3452_ _2740_ _0380_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__nand4_1
XFILLER_0_74_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3934_ _2215_ VGND VGND VPWR VPWR _2226_ sky130_fd_sc_hd__buf_2
XFILLER_0_59_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6722_ _2119_ _1958_ _2280_ _3596_ VGND VGND VPWR VPWR _2283_ sky130_fd_sc_hd__a31o_1
XFILLER_0_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3865_ net194 net33 net44 net26 VGND VGND VPWR VPWR _1471_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6653_ _2445_ _1007_ VGND VGND VPWR VPWR _2207_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5604_ _0911_ _1048_ _1058_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3796_ _0401_ _0707_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6584_ _2129_ _1987_ _2130_ VGND VGND VPWR VPWR _2131_ sky130_fd_sc_hd__a21oi_2
X_5535_ _0982_ _0983_ _0801_ _0803_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5466_ _0739_ net41 _0907_ _0908_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4417_ _3520_ _3436_ VGND VGND VPWR VPWR _3521_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7205_ _2809_ _2810_ VGND VGND VPWR VPWR _2811_ sky130_fd_sc_hd__xor2_1
XFILLER_0_100_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5397_ _0558_ _0559_ _0704_ _0690_ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4348_ _3451_ _3452_ _2106_ _2149_ VGND VGND VPWR VPWR _3453_ sky130_fd_sc_hd__nand4_2
X_7136_ _2728_ _2734_ VGND VGND VPWR VPWR _2735_ sky130_fd_sc_hd__xor2_1
X_4279_ _3343_ VGND VGND VPWR VPWR _3385_ sky130_fd_sc_hd__clkbuf_4
X_7067_ _2483_ _2485_ _2659_ VGND VGND VPWR VPWR _2660_ sky130_fd_sc_hd__a21oi_2
X_6018_ _1346_ _1499_ _1510_ VGND VGND VPWR VPWR _1512_ sky130_fd_sc_hd__nand3_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer1 _0526_ VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__buf_1
X_5320_ _3442_ net36 net37 _3635_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__a22o_1
X_5251_ _0671_ _0672_ _0528_ _0530_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4202_ _3307_ _3308_ VGND VGND VPWR VPWR _3309_ sky130_fd_sc_hd__nor2_1
X_5182_ _0594_ _0598_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__xor2_2
XFILLER_0_48_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4133_ net55 _0074_ VGND VGND VPWR VPWR _3241_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4064_ net1 net60 VGND VGND VPWR VPWR _3173_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4966_ _3196_ _3271_ _3644_ _0247_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__nand4_2
XFILLER_0_74_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6705_ _3209_ _2263_ VGND VGND VPWR VPWR _2264_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4897_ _0079_ _0168_ _0169_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__o21bai_1
X_3917_ _2007_ _2018_ _2029_ VGND VGND VPWR VPWR _2040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3848_ _1275_ _0499_ _0401_ _0739_ VGND VGND VPWR VPWR _1286_ sky130_fd_sc_hd__and4_1
X_6636_ _2185_ _2186_ _2043_ _2167_ VGND VGND VPWR VPWR _2188_ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3779_ _0521_ _0445_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__and2b_1
XFILLER_0_15_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6567_ _0419_ _1957_ _1958_ _1962_ _2112_ VGND VGND VPWR VPWR _2113_ sky130_fd_sc_hd__a311o_1
XFILLER_0_132_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5518_ _0963_ _0964_ _0965_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__nand3_1
XFILLER_0_89_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6498_ _3424_ _3512_ _2499_ _2532_ VGND VGND VPWR VPWR _2037_ sky130_fd_sc_hd__nand4_1
X_5449_ _0428_ _1734_ _0571_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__o21a_1
XFILLER_0_100_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7119_ _0063_ _1799_ net20 _0183_ VGND VGND VPWR VPWR _2716_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_57_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_450 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_667 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4820_ _0007_ _0190_ _0198_ _0203_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__a211o_1
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4751_ _0123_ _0127_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__xnor2_1
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4682_ _3650_ _3652_ _3653_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__a21bo_1
X_7470_ _3096_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__buf_2
XFILLER_0_50_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6421_ _1950_ _1951_ VGND VGND VPWR VPWR _1953_ sky130_fd_sc_hd__or2_2
XFILLER_0_153_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6352_ _3430_ _2532_ _1874_ _1875_ VGND VGND VPWR VPWR _1878_ sky130_fd_sc_hd__o2bb2a_1
X_5303_ _0725_ _0729_ _0730_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__or3_1
X_6283_ _1796_ _1801_ VGND VGND VPWR VPWR _1802_ sky130_fd_sc_hd__nand2_1
X_5234_ _0324_ net163 _0452_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__and3_1
X_5165_ _0560_ _0580_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__nor2_1
X_4116_ _1832_ _2040_ _0947_ VGND VGND VPWR VPWR _3224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5096_ _0503_ _0504_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__nor2_1
X_4047_ _0838_ _1701_ VGND VGND VPWR VPWR _3156_ sky130_fd_sc_hd__nand2_4
XFILLER_0_148_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5998_ _2313_ _0720_ _0873_ _0095_ VGND VGND VPWR VPWR _1490_ sky130_fd_sc_hd__a22o_1
X_4949_ _0342_ _0343_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__or2_4
XFILLER_0_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6619_ _2013_ _2021_ VGND VGND VPWR VPWR _2169_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap107 _1191_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__buf_1
XFILLER_0_52_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap118 _1088_ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__buf_1
XFILLER_0_123_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6970_ _2550_ _2551_ _2552_ VGND VGND VPWR VPWR _2553_ sky130_fd_sc_hd__nand3_4
X_5921_ _1233_ _1235_ _1234_ VGND VGND VPWR VPWR _1407_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5852_ _1330_ VGND VGND VPWR VPWR _1331_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4803_ _3722_ _3724_ _0177_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__o21bai_1
X_5783_ net107 _1192_ _1254_ _1255_ VGND VGND VPWR VPWR _1256_ sky130_fd_sc_hd__or4_4
XFILLER_0_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4734_ net35 VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4665_ _2368_ _3433_ _3431_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__and3_1
X_7453_ _0696_ _0309_ _3075_ _0641_ VGND VGND VPWR VPWR _3080_ sky130_fd_sc_hd__o22a_1
X_7384_ _3001_ _3005_ VGND VGND VPWR VPWR _3006_ sky130_fd_sc_hd__xnor2_1
X_4596_ _3108_ _3698_ VGND VGND VPWR VPWR _3699_ sky130_fd_sc_hd__or2_2
XFILLER_0_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6404_ _1608_ _1756_ VGND VGND VPWR VPWR _1935_ sky130_fd_sc_hd__and2b_1
XFILLER_0_141_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6335_ _1856_ _1857_ _1858_ VGND VGND VPWR VPWR _1859_ sky130_fd_sc_hd__nand3_1
XFILLER_0_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6266_ _1770_ _1782_ _1783_ VGND VGND VPWR VPWR _1784_ sky130_fd_sc_hd__o21a_1
X_5217_ _0633_ _0634_ _0635_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__a21o_1
X_6197_ _1705_ _1706_ _1707_ VGND VGND VPWR VPWR _1708_ sky130_fd_sc_hd__nand3_1
XFILLER_0_98_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5148_ _0560_ _0561_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__or2_1
X_5079_ _0465_ _0467_ _0484_ _0485_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_67_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_751 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4450_ _3519_ _3552_ _3553_ VGND VGND VPWR VPWR _3554_ sky130_fd_sc_hd__and3_4
XFILLER_0_123_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4381_ _3108_ VGND VGND VPWR VPWR _3486_ sky130_fd_sc_hd__clkbuf_4
X_6120_ _1601_ _1599_ _1621_ _1622_ VGND VGND VPWR VPWR _1623_ sky130_fd_sc_hd__o211a_2
XFILLER_0_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6051_ _3631_ _2773_ _1546_ _1547_ VGND VGND VPWR VPWR _1549_ sky130_fd_sc_hd__nand4_1
XFILLER_0_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _0331_ _0400_ _0402_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__or3_4
XFILLER_0_56_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6953_ _2522_ _2523_ _2533_ VGND VGND VPWR VPWR _2535_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_72_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5904_ _3633_ net7 net8 _3195_ VGND VGND VPWR VPWR _1388_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6884_ _0357_ _1949_ _2458_ _2459_ VGND VGND VPWR VPWR _2460_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_76_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5835_ _3589_ _1297_ _1277_ VGND VGND VPWR VPWR _1312_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_146_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5766_ _1234_ _1235_ _1233_ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4717_ _0018_ _0027_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__and2b_1
XFILLER_0_115_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5697_ _1160_ VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4648_ net138 VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7436_ _3587_ _3050_ _3051_ _3054_ _3061_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__a2111o_4
XFILLER_0_16_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4579_ _3610_ _3681_ VGND VGND VPWR VPWR _3682_ sky130_fd_sc_hd__xor2_1
X_7367_ _2983_ _2986_ VGND VGND VPWR VPWR _2987_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7298_ _2909_ _2910_ VGND VGND VPWR VPWR _2911_ sky130_fd_sc_hd__nor2_1
X_6318_ _1660_ _1667_ _1666_ VGND VGND VPWR VPWR _1840_ sky130_fd_sc_hd__a21bo_1
X_6249_ _1609_ _1764_ VGND VGND VPWR VPWR _1765_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_843 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3950_ _2390_ VGND VGND VPWR VPWR _2401_ sky130_fd_sc_hd__buf_4
XFILLER_0_133_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3881_ _1613_ _1635_ VGND VGND VPWR VPWR _1646_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5620_ _1075_ _1076_ VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5551_ _0878_ _1001_ _0181_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4502_ _3596_ _3600_ _3601_ _3605_ _0860_ VGND VGND VPWR VPWR _3606_ sky130_fd_sc_hd__o32a_1
XFILLER_0_13_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5482_ _0769_ _0777_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__nand2_1
X_7221_ _2335_ _2401_ _1607_ _1797_ VGND VGND VPWR VPWR _2829_ sky130_fd_sc_hd__and4_1
XFILLER_0_41_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4433_ net2 VGND VGND VPWR VPWR _3537_ sky130_fd_sc_hd__buf_4
XFILLER_0_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4364_ _3466_ _3467_ _3427_ VGND VGND VPWR VPWR _3469_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7152_ _3685_ _2609_ VGND VGND VPWR VPWR _2753_ sky130_fd_sc_hd__nand2_1
X_4295_ _1985_ _2631_ _1712_ VGND VGND VPWR VPWR _3401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7083_ _2311_ _2677_ _2672_ VGND VGND VPWR VPWR _2678_ sky130_fd_sc_hd__a21o_1
X_6103_ _1458_ _1459_ _1472_ _1605_ VGND VGND VPWR VPWR _1606_ sky130_fd_sc_hd__a211o_1
X_6034_ _3423_ _0105_ _2696_ _2751_ VGND VGND VPWR VPWR _1530_ sky130_fd_sc_hd__nand4_4
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer11 _0650_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__buf_1
XFILLER_0_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer55 _0405_ VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_1
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer22 _3257_ VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer33 _2098_ VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__buf_1
Xrebuffer44 _2493_ VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer66 _0267_ VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_692 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6936_ _2903_ _1745_ VGND VGND VPWR VPWR _2516_ sky130_fd_sc_hd__nand2_1
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer77 _2397_ VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6867_ _2397_ _2398_ _2438_ _2439_ VGND VGND VPWR VPWR _2441_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_9_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5818_ _1268_ _1269_ _1293_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__o21ai_4
X_6798_ _2355_ _2364_ VGND VGND VPWR VPWR _2365_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5749_ _0042_ _2773_ _1103_ _1102_ _2532_ VGND VGND VPWR VPWR _1218_ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7419_ _2900_ _3042_ _3043_ VGND VGND VPWR VPWR _3044_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_802 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput91 net91 VGND VGND VPWR VPWR result[2] sky130_fd_sc_hd__clkbuf_4
Xoutput80 net80 VGND VGND VPWR VPWR result[1] sky130_fd_sc_hd__clkbuf_4
X_4080_ _1439_ _3188_ VGND VGND VPWR VPWR _3189_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4982_ _3448_ _2740_ _0380_ _3449_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3933_ _2204_ VGND VGND VPWR VPWR _2215_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6721_ _2119_ _1958_ _2280_ VGND VGND VPWR VPWR _2282_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_144_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3864_ net194 net26 net33 net44 VGND VGND VPWR VPWR _1460_ sky130_fd_sc_hd__and4_1
XFILLER_0_6_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6652_ _2203_ _2205_ VGND VGND VPWR VPWR _2206_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5603_ _0911_ _1048_ _1058_ VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3795_ _0423_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__buf_4
XFILLER_0_73_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6583_ _1968_ _1984_ VGND VGND VPWR VPWR _2130_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5534_ _0801_ _0803_ _0982_ _0983_ VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5465_ _0085_ _1264_ net39 net40 VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__and4_1
XFILLER_0_14_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4416_ _0205_ _0335_ _3196_ _3272_ VGND VGND VPWR VPWR _3520_ sky130_fd_sc_hd__and4_1
XFILLER_0_68_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7204_ _1056_ net54 VGND VGND VPWR VPWR _2810_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7135_ _2730_ _2733_ VGND VGND VPWR VPWR _2734_ sky130_fd_sc_hd__xnor2_1
X_5396_ _0829_ _0831_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__and2_1
X_4347_ _3176_ VGND VGND VPWR VPWR _3452_ sky130_fd_sc_hd__buf_6
X_4278_ _3262_ _3336_ _3381_ _3382_ VGND VGND VPWR VPWR _3384_ sky130_fd_sc_hd__or4bb_4
X_7066_ _2657_ _2658_ VGND VGND VPWR VPWR _2659_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6017_ _1346_ _1499_ _1510_ VGND VGND VPWR VPWR _1511_ sky130_fd_sc_hd__a21o_1
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6919_ _0320_ _2496_ _2497_ VGND VGND VPWR VPWR _2498_ sky130_fd_sc_hd__and3_1
XFILLER_0_147_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer2 _3682_ VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5250_ _0528_ _0530_ _0671_ _0672_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__a211oi_2
X_4201_ net163 net1 _3196_ _3271_ VGND VGND VPWR VPWR _3308_ sky130_fd_sc_hd__and4_1
X_5181_ _3719_ _0595_ _0596_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_48_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4132_ _3238_ _3239_ VGND VGND VPWR VPWR _3240_ sky130_fd_sc_hd__xnor2_2
X_4063_ _3170_ _3171_ VGND VGND VPWR VPWR _3172_ sky130_fd_sc_hd__nor2_2
XFILLER_0_64_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4965_ _3271_ _2106_ _2149_ _3632_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3916_ _0881_ VGND VGND VPWR VPWR _2029_ sky130_fd_sc_hd__buf_6
X_6704_ net52 VGND VGND VPWR VPWR _2263_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4896_ _0286_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6635_ _2043_ _2167_ _2185_ net117 VGND VGND VPWR VPWR _2187_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_62_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3847_ _1264_ VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__buf_4
XFILLER_0_15_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3778_ _0401_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6566_ _2110_ _2111_ _0320_ VGND VGND VPWR VPWR _2112_ sky130_fd_sc_hd__and3b_1
XFILLER_0_131_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5517_ _3451_ _3448_ _2565_ _2598_ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__nand4_2
XFILLER_0_14_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6497_ _2034_ _2035_ VGND VGND VPWR VPWR _2036_ sky130_fd_sc_hd__xor2_2
XFILLER_0_30_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5448_ _0855_ _0876_ _0877_ _0854_ _0888_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5379_ _0673_ _0718_ _0812_ _0813_ VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__o211a_2
X_7118_ _2711_ _2712_ _2713_ VGND VGND VPWR VPWR _2715_ sky130_fd_sc_hd__a21o_1
X_7049_ _2462_ _2627_ _2638_ _2639_ VGND VGND VPWR VPWR _2640_ sky130_fd_sc_hd__a211oi_4
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_495 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _0124_ _0126_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__xor2_2
XFILLER_0_56_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4681_ _0049_ _0050_ _0048_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6420_ _1810_ _1949_ VGND VGND VPWR VPWR _1951_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6351_ _1874_ _1875_ _3343_ _2521_ VGND VGND VPWR VPWR _1877_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_12_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5302_ _0423_ _0654_ _0726_ _0727_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_52_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6282_ _1798_ _1800_ VGND VGND VPWR VPWR _1801_ sky130_fd_sc_hd__nor2_1
X_5233_ _0466_ _0654_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__nand2_1
X_5164_ _0438_ _0579_ _0000_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__a21oi_1
X_4115_ _3219_ _3220_ _3221_ _3222_ _1712_ _1723_ VGND VGND VPWR VPWR _3223_ sky130_fd_sc_hd__mux4_1
X_5095_ _3645_ _0041_ _0491_ _2686_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__and4_1
X_4046_ _3108_ _3145_ _3153_ _1734_ _3154_ VGND VGND VPWR VPWR _3155_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5997_ _0095_ _2313_ _0720_ _0873_ VGND VGND VPWR VPWR _1489_ sky130_fd_sc_hd__and4_1
XFILLER_0_148_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4948_ _0338_ _0341_ _0434_ _0219_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4879_ _0246_ _0266_ _0267_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6618_ _2020_ _2014_ VGND VGND VPWR VPWR _2168_ sky130_fd_sc_hd__and2b_1
XFILLER_0_46_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6549_ _1910_ net103 _2091_ _2092_ VGND VGND VPWR VPWR _2093_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap108 _1737_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__buf_2
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap119 _0979_ VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5920_ _1401_ _1402_ _1403_ VGND VGND VPWR VPWR _1405_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5851_ _0085_ _1264_ net42 net43 VGND VGND VPWR VPWR _1330_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4802_ _3722_ _3724_ _0177_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__or3b_1
X_5782_ _1251_ _1252_ _1124_ net137 VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4733_ _0107_ _0108_ _0739_ _3619_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_28_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7452_ _3078_ VGND VGND VPWR VPWR _3079_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4664_ _0095_ _3631_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6403_ _1932_ _1933_ VGND VGND VPWR VPWR _1934_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7383_ _3003_ _3004_ VGND VGND VPWR VPWR _3005_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4595_ _0554_ _3291_ _3035_ _3144_ VGND VGND VPWR VPWR _3698_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_43_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6334_ _1703_ _1704_ _1702_ VGND VGND VPWR VPWR _1858_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_101_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6265_ _1770_ _1782_ _0181_ VGND VGND VPWR VPWR _1783_ sky130_fd_sc_hd__a21oi_1
X_5216_ _0633_ _0634_ _0635_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__nand3_2
XFILLER_0_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6196_ _1556_ _1557_ _1555_ VGND VGND VPWR VPWR _1707_ sky130_fd_sc_hd__a21bo_1
X_5147_ _0558_ _0559_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__and2_1
X_5078_ _0482_ _0483_ _0468_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__a21oi_1
X_4029_ _2182_ _2237_ _3137_ _2675_ _0914_ _0958_ VGND VGND VPWR VPWR _3138_ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsplit38 _3270_ VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__buf_2
XFILLER_0_149_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4380_ _3482_ _3483_ VGND VGND VPWR VPWR _3485_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6050_ _3633_ net8 _2521_ _3195_ VGND VGND VPWR VPWR _1547_ sky130_fd_sc_hd__a22o_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ net115 _0399_ net156 _0273_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6952_ _2522_ _2523_ _2533_ VGND VGND VPWR VPWR _2534_ sky130_fd_sc_hd__or3_1
X_5903_ _3632_ _3633_ _0380_ _2489_ VGND VGND VPWR VPWR _1387_ sky130_fd_sc_hd__nand4_2
XFILLER_0_72_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6883_ _0106_ _0215_ _1607_ net50 VGND VGND VPWR VPWR _2459_ sky130_fd_sc_hd__and4_1
XFILLER_0_146_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5834_ _0844_ _1310_ _3228_ VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_146_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5765_ _1233_ _1234_ _1235_ VGND VGND VPWR VPWR _1236_ sky130_fd_sc_hd__nand3_1
XFILLER_0_44_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4716_ _3612_ net149 _3675_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__nand3_1
XFILLER_0_115_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5696_ _1264_ _0314_ net42 net43 VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__and4_1
XFILLER_0_8_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4647_ _0015_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7435_ _3055_ _2980_ _3057_ _3060_ VGND VGND VPWR VPWR _3061_ sky130_fd_sc_hd__a31o_1
XFILLER_0_71_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7366_ _2984_ _2985_ VGND VGND VPWR VPWR _2986_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4578_ _3679_ _3680_ VGND VGND VPWR VPWR _3681_ sky130_fd_sc_hd__nand2_2
X_6317_ _1836_ _1837_ _1830_ VGND VGND VPWR VPWR _1839_ sky130_fd_sc_hd__a21o_1
X_7297_ _2758_ _2908_ _3137_ _1008_ VGND VGND VPWR VPWR _2910_ sky130_fd_sc_hd__o211a_1
X_6248_ _0438_ _1763_ _0000_ VGND VGND VPWR VPWR _1764_ sky130_fd_sc_hd__a21oi_1
X_6179_ _3511_ _2740_ _0380_ _3422_ VGND VGND VPWR VPWR _1688_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3880_ _1406_ _1624_ VGND VGND VPWR VPWR _1635_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5550_ _0829_ _0831_ _1000_ VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5481_ _0770_ _0774_ _0775_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__or3_1
X_4501_ _1734_ _3604_ VGND VGND VPWR VPWR _3605_ sky130_fd_sc_hd__or2b_1
XFILLER_0_130_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4432_ _0292_ _2106_ VGND VGND VPWR VPWR _3536_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7220_ _2401_ _1608_ _1797_ _2335_ VGND VGND VPWR VPWR _2827_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_111_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4363_ _3427_ _3466_ _3467_ VGND VGND VPWR VPWR _3468_ sky130_fd_sc_hd__nand3_2
X_7151_ _2749_ _2750_ VGND VGND VPWR VPWR _2752_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6102_ _0320_ _1602_ _1604_ VGND VGND VPWR VPWR _1605_ sky130_fd_sc_hd__and3_1
X_4294_ _2292_ _2806_ _1100_ VGND VGND VPWR VPWR _3400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7082_ _2299_ _2007_ VGND VGND VPWR VPWR _2677_ sky130_fd_sc_hd__or2b_1
X_6033_ _3424_ _3512_ _2653_ _2707_ VGND VGND VPWR VPWR _1529_ sky130_fd_sc_hd__and4_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer12 _1126_ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__buf_1
Xrebuffer23 _3257_ VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer34 _2098_ VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_1
Xrebuffer45 _2096_ VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__buf_1
Xrebuffer56 net181 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6935_ _2513_ _2514_ VGND VGND VPWR VPWR _2515_ sky130_fd_sc_hd__nor2_1
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer67 _1121_ VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_1
Xrebuffer78 _1251_ VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__buf_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6866_ _2397_ _2398_ _2438_ _2439_ VGND VGND VPWR VPWR _2440_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_147_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6797_ _2362_ _2363_ VGND VGND VPWR VPWR _2364_ sky130_fd_sc_hd__and2b_1
X_5817_ _3571_ _1276_ _1292_ VGND VGND VPWR VPWR _1293_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5748_ _3197_ _3272_ _2707_ _2751_ _1097_ VGND VGND VPWR VPWR _1217_ sky130_fd_sc_hd__a41o_1
XFILLER_0_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5679_ _1140_ _1141_ VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7418_ _2900_ _3042_ _3192_ VGND VGND VPWR VPWR _3043_ sky130_fd_sc_hd__a21oi_1
X_7349_ _2965_ _2966_ VGND VGND VPWR VPWR _2967_ sky130_fd_sc_hd__xnor2_1
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_814 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput70 net70 VGND VGND VPWR VPWR result[10] sky130_fd_sc_hd__clkbuf_4
Xoutput92 net92 VGND VGND VPWR VPWR result[30] sky130_fd_sc_hd__buf_2
Xoutput81 net81 VGND VGND VPWR VPWR result[20] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4981_ net7 VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3932_ net2 VGND VGND VPWR VPWR _2204_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6720_ _2278_ _2279_ VGND VGND VPWR VPWR _2280_ sky130_fd_sc_hd__nand2_2
XFILLER_0_144_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3863_ _0303_ _0434_ _1296_ _1286_ VGND VGND VPWR VPWR _1449_ sky130_fd_sc_hd__a31o_1
XFILLER_0_74_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6651_ _2160_ _0721_ _0874_ _2117_ VGND VGND VPWR VPWR _2205_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5602_ _1049_ _1057_ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6582_ _1968_ _1984_ VGND VGND VPWR VPWR _2129_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5533_ _0944_ _0945_ _0979_ _0981_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__o22ai_2
X_3794_ _0499_ _0477_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__nand2_2
XFILLER_0_6_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5464_ _0085_ _0325_ _0452_ _0194_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__a22oi_1
X_4415_ _3517_ _3518_ VGND VGND VPWR VPWR _3519_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5395_ _0829_ _0831_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__nor2_1
X_7203_ _2807_ _2808_ VGND VGND VPWR VPWR _2809_ sky130_fd_sc_hd__nor2_1
X_4346_ _3242_ VGND VGND VPWR VPWR _3451_ sky130_fd_sc_hd__buf_6
XFILLER_0_100_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7134_ _2731_ _2732_ VGND VGND VPWR VPWR _2733_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4277_ _3381_ _3382_ _3338_ VGND VGND VPWR VPWR _3383_ sky130_fd_sc_hd__a21bo_1
X_7065_ _2654_ _2655_ _2656_ VGND VGND VPWR VPWR _2658_ sky130_fd_sc_hd__o21ba_1
X_6016_ _1500_ _1509_ VGND VGND VPWR VPWR _1510_ sky130_fd_sc_hd__xnor2_1
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6918_ net168 _2494_ _2495_ _2491_ VGND VGND VPWR VPWR _2497_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_108_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6849_ _2219_ _2221_ VGND VGND VPWR VPWR _2421_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_560 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer3 net126 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4200_ _0434_ _3196_ _3272_ net1 VGND VGND VPWR VPWR _3307_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_139_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5180_ _3635_ net36 _0340_ _3440_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__a22o_1
X_4131_ _0412_ net60 VGND VGND VPWR VPWR _3239_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4062_ net58 net59 net23 net12 VGND VGND VPWR VPWR _3171_ sky130_fd_sc_hd__and4_1
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4964_ _0249_ _0250_ _0251_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_93_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6703_ _2258_ _2261_ VGND VGND VPWR VPWR _2262_ sky130_fd_sc_hd__xor2_1
X_3915_ net22 VGND VGND VPWR VPWR _2018_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_129_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4895_ _0207_ _0285_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3846_ net26 VGND VGND VPWR VPWR _1264_ sky130_fd_sc_hd__buf_4
X_6634_ _2168_ _2169_ _2184_ VGND VGND VPWR VPWR _2186_ sky130_fd_sc_hd__nor3_1
XFILLER_0_61_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3777_ _0477_ _0499_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__or2b_2
XFILLER_0_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6565_ _2107_ _2109_ _2105_ VGND VGND VPWR VPWR _2111_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5516_ _0390_ net10 net11 _0488_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__a22o_1
X_6496_ _0178_ _0337_ VGND VGND VPWR VPWR _2035_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_451 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5447_ _0578_ _0885_ _0886_ _0887_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5378_ _0810_ _0811_ _0719_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4329_ _0194_ _0314_ _3433_ _3431_ VGND VGND VPWR VPWR _3434_ sky130_fd_sc_hd__nand4_1
X_7117_ _2711_ _2712_ _2713_ VGND VGND VPWR VPWR _2714_ sky130_fd_sc_hd__nand3_1
X_7048_ _2413_ _2416_ _2637_ VGND VGND VPWR VPWR _2639_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4680_ _0048_ _0049_ _0050_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__nand3_1
XFILLER_0_153_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6350_ _3633_ net10 net11 _3195_ VGND VGND VPWR VPWR _1875_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_52_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5301_ _0726_ _0727_ _0423_ net41 VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_12_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6281_ _0445_ _0991_ _1607_ net50 VGND VGND VPWR VPWR _1800_ sky130_fd_sc_hd__and4_1
XFILLER_0_121_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5232_ net41 VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__buf_2
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5163_ _0558_ _0559_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__nand2_1
X_4114_ _2467_ _2193_ _3131_ VGND VGND VPWR VPWR _3222_ sky130_fd_sc_hd__mux2_1
X_5094_ _0041_ _0491_ _2696_ _3645_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__a22oi_2
X_4045_ _1154_ _1144_ _1165_ VGND VGND VPWR VPWR _3154_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_79_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5996_ _1485_ _1487_ VGND VGND VPWR VPWR _1488_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4947_ _1428_ _0337_ _0338_ _0341_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4878_ _0263_ _0264_ _0265_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6617_ _2036_ _2045_ VGND VGND VPWR VPWR _2167_ sky130_fd_sc_hd__or2_1
X_3829_ _1023_ _1034_ _1045_ _1067_ _0903_ _0947_ VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__mux4_1
XFILLER_0_7_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6548_ _2054_ _2055_ _2089_ _2090_ VGND VGND VPWR VPWR _2092_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_42_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6479_ _3272_ _2598_ _1854_ _3196_ VGND VGND VPWR VPWR _2016_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_30_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_579 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap109 _1420_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__buf_1
XFILLER_0_104_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap1 _2849_ VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5850_ _1326_ _1327_ VGND VGND VPWR VPWR _1328_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4801_ _0177_ _0180_ _0182_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__o21a_1
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5781_ _1124_ net137 net214 _1252_ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_28_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4732_ _0085_ _0194_ _3422_ _3511_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__and4_1
XFILLER_0_84_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4663_ _3643_ _3646_ _3647_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__o21ba_1
X_7451_ _0863_ _3209_ _0855_ _3076_ _1277_ VGND VGND VPWR VPWR _3078_ sky130_fd_sc_hd__o32a_1
XFILLER_0_43_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6402_ _1763_ _1615_ _1930_ _3596_ VGND VGND VPWR VPWR _1933_ sky130_fd_sc_hd__a31o_1
X_7382_ _3513_ _1909_ VGND VGND VPWR VPWR _3004_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4594_ _3296_ _3299_ _3292_ _3298_ _3301_ _3490_ VGND VGND VPWR VPWR _3697_ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6333_ _1852_ _1853_ _1855_ VGND VGND VPWR VPWR _1857_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6264_ _0567_ _1771_ _1772_ _1781_ VGND VGND VPWR VPWR _1782_ sky130_fd_sc_hd__a31o_1
X_5215_ _0507_ _0508_ _0509_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_86_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6195_ _1702_ _1703_ _1704_ VGND VGND VPWR VPWR _1706_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5146_ _0558_ _0559_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__nor2_1
X_5077_ _0468_ _0482_ _0483_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4028_ _2270_ VGND VGND VPWR VPWR _3137_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsplit39 _0412_ VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_2
X_5979_ _0844_ _1468_ VGND VGND VPWR VPWR _1469_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5000_ net156 _0273_ net172 _0399_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__a211oi_4
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6951_ _2524_ _2531_ VGND VGND VPWR VPWR _2533_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5902_ _2881_ _2489_ _1228_ _1227_ _2565_ VGND VGND VPWR VPWR _1386_ sky130_fd_sc_hd__a32o_1
XFILLER_0_72_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6882_ _0106_ _1607_ net50 _0215_ VGND VGND VPWR VPWR _2458_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_146_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5833_ _0305_ _1309_ _0867_ VGND VGND VPWR VPWR _1310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5764_ _0390_ net13 _1887_ _0488_ VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4715_ _0089_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_6
XFILLER_0_71_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5695_ _1059_ _1061_ VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__nor2_1
X_4646_ _3626_ _3615_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__and2b_1
XFILLER_0_115_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7434_ _0685_ _3058_ _3059_ _0652_ VGND VGND VPWR VPWR _3060_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4577_ _3676_ _3677_ _3678_ VGND VGND VPWR VPWR _3680_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7365_ _2777_ _2778_ _2776_ VGND VGND VPWR VPWR _2985_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_13_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6316_ _1830_ _1836_ _1837_ VGND VGND VPWR VPWR _1838_ sky130_fd_sc_hd__nand3_2
XFILLER_0_110_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7296_ _3137_ _1008_ _2758_ _2908_ VGND VGND VPWR VPWR _2909_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_40_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6247_ _1756_ _1608_ VGND VGND VPWR VPWR _1763_ sky130_fd_sc_hd__nand2_1
X_6178_ _0104_ _3511_ _2740_ _0380_ VGND VGND VPWR VPWR _1687_ sky130_fd_sc_hd__nand4_2
X_5129_ _0538_ _0539_ _0446_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5480_ _0754_ _0762_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__and2_2
XFILLER_0_81_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4500_ _3212_ _3603_ _3301_ VGND VGND VPWR VPWR _3604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4431_ _2925_ _3534_ VGND VGND VPWR VPWR _3535_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_1 _1753_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4362_ _3464_ _3465_ _3368_ net122 VGND VGND VPWR VPWR _3467_ sky130_fd_sc_hd__a211o_1
X_7150_ _3425_ _3513_ _1865_ _1898_ VGND VGND VPWR VPWR _2750_ sky130_fd_sc_hd__and4_1
XFILLER_0_67_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4293_ _3389_ _3397_ _2980_ VGND VGND VPWR VPWR _3399_ sky130_fd_sc_hd__o21a_1
X_6101_ _1444_ _1601_ _1599_ _1600_ VGND VGND VPWR VPWR _1604_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7081_ _2672_ _2673_ _2674_ VGND VGND VPWR VPWR _2676_ sky130_fd_sc_hd__o21a_1
X_6032_ _1525_ _1527_ VGND VGND VPWR VPWR _1528_ sky130_fd_sc_hd__xor2_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer24 _3674_ VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_1
Xrebuffer35 _3255_ VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__buf_1
Xrebuffer13 _1126_ VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__buf_6
Xrebuffer46 _2096_ VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_1
Xrebuffer57 _0408_ VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_1
Xrebuffer68 _3334_ VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__buf_1
XFILLER_0_107_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer79 net106 VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__dlymetal6s2s_1
X_6934_ _0172_ _0052_ _1767_ _1799_ VGND VGND VPWR VPWR _2514_ sky130_fd_sc_hd__and4_1
XFILLER_0_49_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6865_ _2436_ _2437_ _2399_ _2229_ VGND VGND VPWR VPWR _2439_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6796_ _2360_ _2361_ _2356_ VGND VGND VPWR VPWR _2363_ sky130_fd_sc_hd__a21o_1
X_5816_ _1282_ _1288_ _1291_ VGND VGND VPWR VPWR _1292_ sky130_fd_sc_hd__or3b_2
XFILLER_0_146_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5747_ _1213_ _1214_ _1193_ _1194_ VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5678_ _0814_ _0994_ _0993_ VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__a21oi_1
X_7417_ _3023_ _3041_ VGND VGND VPWR VPWR _3042_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4629_ _3727_ _3730_ VGND VGND VPWR VPWR _3731_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7348_ _2138_ _1448_ VGND VGND VPWR VPWR _2966_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7279_ _0571_ _2018_ _2051_ _2007_ _0864_ _0863_ VGND VGND VPWR VPWR _2890_ sky130_fd_sc_hd__mux4_1
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput82 net82 VGND VGND VPWR VPWR result[21] sky130_fd_sc_hd__clkbuf_4
Xoutput71 net71 VGND VGND VPWR VPWR result[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput93 net93 VGND VGND VPWR VPWR result[31] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4980_ _0292_ _2686_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3931_ _2138_ _2182_ _2029_ VGND VGND VPWR VPWR _2193_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3862_ _0587_ _0827_ _1428_ _0466_ VGND VGND VPWR VPWR _1439_ sky130_fd_sc_hd__or4b_4
XFILLER_0_86_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6650_ _2117_ _2160_ _0721_ _0874_ VGND VGND VPWR VPWR _2203_ sky130_fd_sc_hd__nand4_1
XFILLER_0_144_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5601_ _1054_ _1055_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6581_ net158 _2100_ VGND VGND VPWR VPWR _2128_ sky130_fd_sc_hd__nand2_2
XFILLER_0_144_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5532_ _0944_ _0945_ _0979_ _0981_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__or4_4
X_3793_ _0521_ _0445_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5463_ _0727_ _0729_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4414_ _3509_ _3510_ _3516_ VGND VGND VPWR VPWR _3518_ sky130_fd_sc_hd__or3_1
XFILLER_0_78_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5394_ _0693_ _0695_ _0830_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__a21o_1
X_7202_ _0226_ _1045_ net52 _2299_ VGND VGND VPWR VPWR _2808_ sky130_fd_sc_hd__and4_1
XFILLER_0_41_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4345_ _3448_ net31 net32 _3449_ VGND VGND VPWR VPWR _3450_ sky130_fd_sc_hd__a22o_1
X_7133_ _3198_ _3273_ _1952_ _1745_ VGND VGND VPWR VPWR _2732_ sky130_fd_sc_hd__and4_1
XFILLER_0_78_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4276_ _3259_ net192 net188 _3380_ VGND VGND VPWR VPWR _3382_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_94_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7064_ _2654_ _2655_ _2656_ VGND VGND VPWR VPWR _2657_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_94_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6015_ _1507_ _1508_ VGND VGND VPWR VPWR _1509_ sky130_fd_sc_hd__and2b_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6917_ _2491_ _2493_ _2494_ _2495_ VGND VGND VPWR VPWR _2496_ sky130_fd_sc_hd__or4_1
XFILLER_0_147_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6848_ _2217_ _2224_ VGND VGND VPWR VPWR _2420_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6779_ _0052_ _1745_ _1767_ _0183_ VGND VGND VPWR VPWR _2344_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_45_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_699 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer4 net207 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__buf_1
XFILLER_0_3_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4130_ _3236_ _3237_ VGND VGND VPWR VPWR _3238_ sky130_fd_sc_hd__nor2_1
X_4061_ _3169_ _0314_ _0412_ net191 VGND VGND VPWR VPWR _3170_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4963_ _2390_ _3385_ _0242_ _0241_ _3197_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__a32o_1
XFILLER_0_74_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3914_ net21 VGND VGND VPWR VPWR _2007_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6702_ _1802_ _1979_ _2260_ VGND VGND VPWR VPWR _2261_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_46_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4894_ _0282_ _0284_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6633_ _2168_ _2169_ _2184_ VGND VGND VPWR VPWR _2185_ sky130_fd_sc_hd__o21a_2
XFILLER_0_144_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3845_ _0128_ _1176_ _1187_ _0139_ _1242_ VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3776_ _0488_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__buf_6
XFILLER_0_70_840 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6564_ _2105_ _2107_ _2109_ VGND VGND VPWR VPWR _2110_ sky130_fd_sc_hd__and3_1
X_5515_ _0281_ _2521_ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__and2_1
X_6495_ _2032_ _2033_ VGND VGND VPWR VPWR _2034_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5446_ _0862_ _0875_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5377_ _0719_ _0810_ _0811_ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7116_ _2504_ _2506_ _2505_ VGND VGND VPWR VPWR _2713_ sky130_fd_sc_hd__a21bo_1
X_4328_ net61 VGND VGND VPWR VPWR _3433_ sky130_fd_sc_hd__clkbuf_4
X_4259_ _3356_ _3363_ _3364_ VGND VGND VPWR VPWR _3365_ sky130_fd_sc_hd__nand3_1
X_7047_ _2413_ _2416_ _2637_ VGND VGND VPWR VPWR _2638_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_69_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5300_ _0194_ _0324_ _0325_ _0452_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__and4_1
XFILLER_0_51_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6280_ _1056_ _1607_ _1797_ _0991_ VGND VGND VPWR VPWR _1798_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_121_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5231_ _0346_ _0220_ _0471_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__and3_1
X_5162_ _0783_ _3156_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__nor2_2
XFILLER_0_20_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5093_ _0042_ _2259_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__nand2_1
X_4113_ _2281_ _2729_ _3131_ VGND VGND VPWR VPWR _3221_ sky130_fd_sc_hd__mux2_1
X_4044_ _0870_ _3152_ VGND VGND VPWR VPWR _3153_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5995_ _0991_ net48 _1483_ _1486_ VGND VGND VPWR VPWR _1487_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_115_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4946_ _1275_ _0739_ _0339_ _0340_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__and4_1
XFILLER_0_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4877_ _0263_ _0264_ _0265_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__nand3_4
XFILLER_0_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6616_ _2163_ _2164_ _2011_ _2132_ VGND VGND VPWR VPWR _2166_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_7_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3828_ _1056_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__buf_4
XFILLER_0_145_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6547_ _2054_ _2055_ _2089_ _2090_ VGND VGND VPWR VPWR _2091_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_132_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3759_ net23 VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__buf_8
XFILLER_0_15_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6478_ _3196_ _3272_ _2598_ _1854_ VGND VGND VPWR VPWR _2015_ sky130_fd_sc_hd__and4_1
XFILLER_0_30_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5429_ _3283_ _3702_ _0433_ _0865_ _0866_ _0867_ VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__mux4_1
XFILLER_0_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap2 _1324_ VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4800_ _0177_ _0180_ _0181_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_145_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5780_ _1215_ _1216_ _1249_ _1250_ VGND VGND VPWR VPWR _1252_ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_0_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4731_ _3440_ _0104_ _0105_ _0194_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_72_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4662_ _3636_ _3637_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__nand2_2
X_7450_ _3305_ _0696_ _0438_ _3075_ VGND VGND VPWR VPWR _3076_ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6401_ _1763_ _1615_ _1930_ VGND VGND VPWR VPWR _1932_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7381_ _3425_ _1942_ VGND VGND VPWR VPWR _3003_ sky130_fd_sc_hd__nand2_1
X_4593_ _3695_ VGND VGND VPWR VPWR _3696_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6332_ _1852_ _1853_ _1855_ VGND VGND VPWR VPWR _1856_ sky130_fd_sc_hd__nand3_1
XFILLER_0_12_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6263_ _1963_ _1773_ _1771_ _1776_ _1780_ VGND VGND VPWR VPWR _1781_ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5214_ _0631_ _0632_ _0629_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6194_ _1702_ _1703_ _1704_ VGND VGND VPWR VPWR _1705_ sky130_fd_sc_hd__nand3_1
XFILLER_0_86_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5145_ _0454_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5076_ _0480_ _0481_ _0473_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4027_ _3133_ _3134_ _3135_ _2510_ _0914_ _0958_ VGND VGND VPWR VPWR _3136_ sky130_fd_sc_hd__mux4_2
XFILLER_0_67_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5978_ _0435_ _1467_ _0867_ VGND VGND VPWR VPWR _1468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4929_ _0232_ _0234_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__or2_2
XFILLER_0_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_618 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_506 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6950_ _2525_ _2530_ VGND VGND VPWR VPWR _2531_ sky130_fd_sc_hd__xor2_2
XFILLER_0_22_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5901_ _1219_ _1222_ VGND VGND VPWR VPWR _1385_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6881_ _2249_ _2251_ VGND VGND VPWR VPWR _2457_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5832_ _0845_ _1308_ _0866_ VGND VGND VPWR VPWR _1309_ sky130_fd_sc_hd__mux2_1
X_5763_ _3451_ _3452_ _1854_ _1887_ VGND VGND VPWR VPWR _1234_ sky130_fd_sc_hd__nand4_2
XFILLER_0_57_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4714_ _3726_ _3732_ _0010_ _0088_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__or4_1
XFILLER_0_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5694_ _1065_ _1066_ _1128_ _1129_ VGND VGND VPWR VPWR _1158_ sky130_fd_sc_hd__nor4_1
XFILLER_0_114_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7433_ _0455_ _0510_ VGND VGND VPWR VPWR _3059_ sky130_fd_sc_hd__xor2_1
X_4645_ _3723_ _0012_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4576_ _3676_ _3677_ _3678_ VGND VGND VPWR VPWR _3679_ sky130_fd_sc_hd__or3_4
XFILLER_0_115_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7364_ _2182_ _1295_ VGND VGND VPWR VPWR _2984_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6315_ _1834_ _1835_ _1683_ _1684_ VGND VGND VPWR VPWR _1837_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_13_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7295_ _2553_ _2556_ _2758_ _2759_ VGND VGND VPWR VPWR _2908_ sky130_fd_sc_hd__a211oi_2
X_6246_ _3156_ _3404_ VGND VGND VPWR VPWR _1762_ sky130_fd_sc_hd__nor2_1
X_6177_ _1684_ _1685_ VGND VGND VPWR VPWR _1686_ sky130_fd_sc_hd__and2_1
X_5128_ _0446_ _0538_ _0539_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__nand3_1
XFILLER_0_99_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5059_ _0449_ _0463_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4430_ _3530_ _3532_ _3533_ VGND VGND VPWR VPWR _3534_ sky130_fd_sc_hd__a21bo_1
XANTENNA_2 _2270_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4361_ _3368_ net122 _3464_ _3465_ VGND VGND VPWR VPWR _3466_ sky130_fd_sc_hd__o211ai_4
X_6100_ _1599_ _1600_ _1444_ _1601_ VGND VGND VPWR VPWR _1602_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_10_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4292_ _3389_ _3397_ VGND VGND VPWR VPWR _3398_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7080_ _2672_ _2673_ _3596_ VGND VGND VPWR VPWR _2674_ sky130_fd_sc_hd__a21oi_1
X_6031_ _2160_ _0220_ VGND VGND VPWR VPWR _1527_ sky130_fd_sc_hd__nand2_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer14 _3666_ VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__buf_1
Xrebuffer25 net148 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__dlygate4sd3_1
Xrebuffer36 net159 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_1
Xrebuffer69 _3233_ VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6933_ _0052_ _1767_ _1799_ _0183_ VGND VGND VPWR VPWR _2513_ sky130_fd_sc_hd__a22oi_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer58 _2094_ VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_1
Xrebuffer47 _2101_ VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__buf_1
X_6864_ _2399_ _2229_ _2436_ _2437_ VGND VGND VPWR VPWR _2438_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_49_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5815_ _1289_ _1290_ VGND VGND VPWR VPWR _1291_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6795_ _2356_ _2360_ _2361_ VGND VGND VPWR VPWR _2362_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5746_ _1193_ _1194_ _1213_ _1214_ VGND VGND VPWR VPWR _1215_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_8_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5677_ _1138_ _1139_ VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4628_ _2073_ _3729_ VGND VGND VPWR VPWR _3730_ sky130_fd_sc_hd__nand2_1
X_7416_ _3025_ _3040_ VGND VGND VPWR VPWR _3041_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4559_ _3659_ _3660_ _3661_ VGND VGND VPWR VPWR _3662_ sky130_fd_sc_hd__nand3_2
X_7347_ _3134_ _0689_ VGND VGND VPWR VPWR _2965_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7278_ _2703_ _2887_ _2883_ VGND VGND VPWR VPWR _2889_ sky130_fd_sc_hd__a21boi_1
X_6229_ _1642_ _1584_ _1741_ _1742_ VGND VGND VPWR VPWR _1743_ sky130_fd_sc_hd__o211ai_2
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput83 net83 VGND VGND VPWR VPWR result[22] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput72 net72 VGND VGND VPWR VPWR result[12] sky130_fd_sc_hd__clkbuf_4
Xoutput94 net94 VGND VGND VPWR VPWR result[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3930_ _2171_ VGND VGND VPWR VPWR _2182_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3861_ _0423_ VGND VGND VPWR VPWR _1428_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3792_ _0183_ _0226_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__nor2_1
X_5600_ _1052_ _1053_ _0929_ _0930_ VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__o211ai_1
X_6580_ _1964_ _2104_ VGND VGND VPWR VPWR _2126_ sky130_fd_sc_hd__nand2_2
XFILLER_0_39_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5531_ _0977_ _0978_ _0797_ _0946_ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5462_ _0901_ _0904_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__and2_1
X_7201_ _0226_ _2263_ _2299_ _1045_ VGND VGND VPWR VPWR _2807_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_112_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4413_ _3509_ _3510_ _3516_ VGND VGND VPWR VPWR _3517_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_78_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5393_ _0689_ _3128_ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4344_ _3242_ VGND VGND VPWR VPWR _3449_ sky130_fd_sc_hd__buf_6
X_7132_ _3273_ _1952_ _1745_ _3198_ VGND VGND VPWR VPWR _2731_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7063_ _2475_ _2479_ VGND VGND VPWR VPWR _2656_ sky130_fd_sc_hd__nand2_1
X_4275_ _3259_ net192 _3379_ _3380_ VGND VGND VPWR VPWR _3381_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_94_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6014_ _1505_ _1506_ _1501_ VGND VGND VPWR VPWR _1508_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6916_ _2102_ _2126_ _2274_ VGND VGND VPWR VPWR _2495_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_147_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6847_ _2218_ _2223_ VGND VGND VPWR VPWR _2419_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6778_ _2339_ _2340_ _2341_ VGND VGND VPWR VPWR _2343_ sky130_fd_sc_hd__a21o_1
XFILLER_0_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5729_ _1092_ _1099_ VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer5 net153 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4060_ net58 VGND VGND VPWR VPWR _3169_ sky130_fd_sc_hd__buf_4
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4962_ _0246_ _0266_ net190 VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__nand3_1
XFILLER_0_129_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4893_ _0073_ _0163_ _0283_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3913_ _1843_ _1985_ _0554_ VGND VGND VPWR VPWR _1996_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6701_ _1978_ _1969_ VGND VGND VPWR VPWR _2260_ sky130_fd_sc_hd__and2b_1
XFILLER_0_144_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3844_ _0139_ _1231_ VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6632_ _2175_ _2183_ VGND VGND VPWR VPWR _2184_ sky130_fd_sc_hd__xor2_1
XFILLER_0_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3775_ net33 VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__clkbuf_4
X_6563_ _1619_ _1620_ _1623_ _2108_ VGND VGND VPWR VPWR _2109_ sky130_fd_sc_hd__a31o_1
XFILLER_0_144_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5514_ _0957_ _0961_ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__xor2_2
XFILLER_0_70_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6494_ _3720_ _2762_ _0191_ VGND VGND VPWR VPWR _2033_ sky130_fd_sc_hd__nand3_1
XFILLER_0_54_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5445_ _3589_ _0877_ _0000_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_14_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5376_ _0808_ _0809_ net135 _0671_ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__a211oi_2
X_7115_ _0980_ net21 _2709_ _2710_ VGND VGND VPWR VPWR _2712_ sky130_fd_sc_hd__nand4_2
X_4327_ _1264_ net61 _3431_ _0314_ VGND VGND VPWR VPWR _3432_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4258_ _3360_ _3361_ _3362_ VGND VGND VPWR VPWR _3364_ sky130_fd_sc_hd__a21o_1
X_7046_ _2628_ _2636_ VGND VGND VPWR VPWR _2637_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4189_ _3130_ _3149_ _0936_ VGND VGND VPWR VPWR _3296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5230_ _0648_ _0649_ _0524_ _0526_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5161_ _0419_ _0569_ _0570_ _0574_ _0575_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__a32o_1
XFILLER_0_20_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5092_ _0490_ _0500_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__xor2_2
X_4112_ _2795_ _2554_ _3131_ VGND VGND VPWR VPWR _3220_ sky130_fd_sc_hd__mux2_1
X_4043_ _3148_ _3151_ _1712_ VGND VGND VPWR VPWR _3152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5994_ _1484_ VGND VGND VPWR VPWR _1486_ sky130_fd_sc_hd__inv_2
X_4945_ net37 VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__buf_4
XFILLER_0_47_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4876_ _0135_ _0144_ _0143_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_74_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6615_ _2011_ _2132_ _2163_ _2164_ VGND VGND VPWR VPWR _2165_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3827_ _0445_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__buf_4
XFILLER_0_131_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3758_ _0292_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__buf_6
XFILLER_0_61_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6546_ _2087_ _2088_ _2056_ VGND VGND VPWR VPWR _2090_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6477_ _2892_ _1865_ _1862_ _1861_ _1931_ VGND VGND VPWR VPWR _2014_ sky130_fd_sc_hd__a32o_1
XFILLER_0_30_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5428_ _0189_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__clkbuf_4
X_5359_ _0788_ _0789_ _0790_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__a21o_1
X_7029_ _1384_ net54 _2616_ _2617_ VGND VGND VPWR VPWR _2618_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_97_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap3 _1158_ VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4730_ _3572_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__buf_4
XFILLER_0_84_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_443 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4661_ _3642_ _3662_ _3663_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__nand3_1
XFILLER_0_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7380_ _0571_ _3046_ VGND VGND VPWR VPWR _3001_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6400_ _1928_ _1929_ VGND VGND VPWR VPWR _1930_ sky130_fd_sc_hd__or2_2
XFILLER_0_43_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6331_ _0292_ net16 VGND VGND VPWR VPWR _1855_ sky130_fd_sc_hd__and2_1
X_4592_ _3573_ _3601_ _3688_ VGND VGND VPWR VPWR _3695_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_12_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6262_ _1452_ _1779_ VGND VGND VPWR VPWR _1780_ sky130_fd_sc_hd__nor2_1
X_5213_ _0629_ _0631_ _0632_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__nand3_1
X_6193_ _0281_ net15 VGND VGND VPWR VPWR _1704_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5144_ _2510_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5075_ _0473_ _0480_ _0481_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__nand3_2
X_4026_ _2784_ VGND VGND VPWR VPWR _3135_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5977_ _0865_ _1466_ _0866_ VGND VGND VPWR VPWR _1467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4928_ _0073_ _0163_ _0282_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__nor3_1
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4859_ _0238_ _0245_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__xor2_2
XFILLER_0_90_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6529_ _1831_ _1834_ VGND VGND VPWR VPWR _2071_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_527 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_616 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5900_ _1226_ _1245_ _1246_ VGND VGND VPWR VPWR _1383_ sky130_fd_sc_hd__nor3_1
XFILLER_0_49_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6880_ _2208_ _2209_ VGND VGND VPWR VPWR _2455_ sky130_fd_sc_hd__or2b_1
X_5831_ _1942_ _1909_ _1876_ _0862_ _0583_ _0864_ VGND VGND VPWR VPWR _1308_ sky130_fd_sc_hd__mux4_1
XFILLER_0_119_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5762_ _0292_ net11 VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4713_ _0652_ _0013_ _0014_ _0087_ _3305_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__a32o_1
XFILLER_0_57_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5693_ _1044_ _1156_ VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_142_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7432_ _0717_ _1209_ _1220_ VGND VGND VPWR VPWR _3058_ sky130_fd_sc_hd__o21ba_1
X_4644_ _3723_ _0012_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4575_ _3473_ _3472_ _3558_ _3559_ VGND VGND VPWR VPWR _3678_ sky130_fd_sc_hd__or4_4
X_7363_ _2725_ _2737_ VGND VGND VPWR VPWR _2983_ sky130_fd_sc_hd__or2b_1
XFILLER_0_12_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7294_ _2901_ _2906_ VGND VGND VPWR VPWR _2907_ sky130_fd_sc_hd__xor2_1
X_6314_ _1683_ _1684_ _1834_ _1835_ VGND VGND VPWR VPWR _1836_ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6245_ _0428_ _1759_ _1760_ _0849_ VGND VGND VPWR VPWR _1761_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6176_ _2215_ _0219_ _1682_ _1683_ VGND VGND VPWR VPWR _1685_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5127_ _0536_ _0537_ _0447_ _0408_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_137_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5058_ _0461_ _0462_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__nand2_1
X_4009_ _0925_ VGND VGND VPWR VPWR _3046_ sky130_fd_sc_hd__buf_4
XFILLER_0_95_814 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_3 _2270_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4360_ _3462_ _3463_ _3439_ VGND VGND VPWR VPWR _3465_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4291_ _3395_ _3396_ VGND VGND VPWR VPWR _3397_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6030_ _3719_ _1523_ _1524_ VGND VGND VPWR VPWR _1525_ sky130_fd_sc_hd__a21bo_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer15 net138 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_1
Xrebuffer26 net148 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer48 net115 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_2
Xrebuffer59 _3372_ VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_1
Xrebuffer37 _1134_ VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_1
X_6932_ _2507_ _2508_ _2509_ VGND VGND VPWR VPWR _2512_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_803 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6863_ _2433_ _2435_ _2185_ _2187_ VGND VGND VPWR VPWR _2437_ sky130_fd_sc_hd__a211o_1
X_5814_ _1021_ _1029_ _1272_ _3596_ VGND VGND VPWR VPWR _1290_ sky130_fd_sc_hd__a31o_1
XFILLER_0_146_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6794_ _3386_ _1865_ _2358_ _2359_ VGND VGND VPWR VPWR _2361_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5745_ _1195_ _1196_ _1212_ VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__nor3_2
XFILLER_0_29_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5676_ _1135_ _1136_ _1137_ VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4627_ _0980_ _0870_ VGND VGND VPWR VPWR _3729_ sky130_fd_sc_hd__nor2_1
X_7415_ _3028_ _3039_ VGND VGND VPWR VPWR _3040_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_698 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4558_ _3535_ _3544_ _3543_ VGND VGND VPWR VPWR _3661_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_114_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7346_ _2957_ _2963_ VGND VGND VPWR VPWR _2964_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4489_ _3574_ _3590_ _3592_ _3201_ VGND VGND VPWR VPWR _3593_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7277_ _2883_ _2887_ _2703_ VGND VGND VPWR VPWR _2888_ sky130_fd_sc_hd__and3b_1
X_6228_ _1678_ _1680_ _1739_ _1740_ VGND VGND VPWR VPWR _1742_ sky130_fd_sc_hd__o22ai_2
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _1661_ _1664_ _1665_ VGND VGND VPWR VPWR _1666_ sky130_fd_sc_hd__nand3_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_646 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput84 net84 VGND VGND VPWR VPWR result[23] sky130_fd_sc_hd__clkbuf_4
Xoutput73 net73 VGND VGND VPWR VPWR result[13] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput95 net165 VGND VGND VPWR VPWR result[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3860_ _0172_ _0707_ _0477_ _0052_ VGND VGND VPWR VPWR _1417_ sky130_fd_sc_hd__a22o_1
X_3791_ _0150_ _0608_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5530_ _0797_ _0946_ _0977_ _0978_ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_82_850 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5461_ _0902_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4412_ _3514_ _3515_ VGND VGND VPWR VPWR _3516_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7200_ _2624_ _2643_ _2644_ VGND VGND VPWR VPWR _2805_ sky130_fd_sc_hd__or3_1
XFILLER_0_42_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5392_ _0826_ _0828_ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__or2_2
XFILLER_0_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4343_ _3176_ VGND VGND VPWR VPWR _3448_ sky130_fd_sc_hd__buf_6
X_7131_ _3386_ _1931_ VGND VGND VPWR VPWR _2730_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4274_ net147 _3334_ _3377_ _3378_ VGND VGND VPWR VPWR _3380_ sky130_fd_sc_hd__o22ai_1
X_7062_ _2651_ _2652_ _2502_ _2481_ VGND VGND VPWR VPWR _2655_ sky130_fd_sc_hd__a211oi_1
X_6013_ _1501_ _1505_ _1506_ VGND VGND VPWR VPWR _1507_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6915_ _2105_ _2107_ _2275_ VGND VGND VPWR VPWR _2494_ sky130_fd_sc_hd__nor3_1
XFILLER_0_76_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_699 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6846_ _2416_ _2417_ VGND VGND VPWR VPWR _2418_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6777_ _2339_ _2340_ _2341_ VGND VGND VPWR VPWR _2342_ sky130_fd_sc_hd__nand3_1
XFILLER_0_91_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3989_ _2095_ _2817_ _0838_ VGND VGND VPWR VPWR _2828_ sky130_fd_sc_hd__mux2_1
X_5728_ _1098_ _1093_ VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__and2b_1
XFILLER_0_60_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5659_ _1116_ _1117_ _1118_ VGND VGND VPWR VPWR _1120_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7329_ _3198_ _1963_ _2944_ VGND VGND VPWR VPWR _2945_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer6 _0984_ VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__buf_1
XFILLER_0_63_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_588 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4961_ _0354_ _0355_ _0332_ _0333_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__o211a_1
X_4892_ _0160_ _0162_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__nand2_1
X_3912_ _1920_ _1974_ _0936_ VGND VGND VPWR VPWR _1985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6700_ _2255_ _2257_ VGND VGND VPWR VPWR _2258_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3843_ _0128_ _1209_ _1220_ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__o21ba_1
X_6631_ _2180_ _2181_ VGND VGND VPWR VPWR _2183_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3774_ _0466_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__buf_4
XFILLER_0_6_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6562_ _1754_ _1926_ VGND VGND VPWR VPWR _2108_ sky130_fd_sc_hd__or2_1
X_5513_ _2489_ _0959_ _0960_ VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_70_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6493_ _3720_ _2751_ _0191_ VGND VGND VPWR VPWR _2032_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5444_ _0884_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__inv_2
X_5375_ net135 _0671_ _0808_ _0809_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__o211a_1
X_7114_ _0980_ net21 _2709_ _2710_ VGND VGND VPWR VPWR _2711_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4326_ _3270_ VGND VGND VPWR VPWR _3431_ sky130_fd_sc_hd__buf_4
XFILLER_0_129_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4257_ _3360_ _3361_ _3362_ VGND VGND VPWR VPWR _3363_ sky130_fd_sc_hd__nand3_1
X_7045_ _2629_ _2635_ VGND VGND VPWR VPWR _2636_ sky130_fd_sc_hd__xnor2_2
X_4188_ _3108_ _3144_ _3200_ _3294_ _3154_ VGND VGND VPWR VPWR _3295_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_145_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6829_ _2214_ _2216_ _2225_ VGND VGND VPWR VPWR _2399_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_37_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_476 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5160_ _0630_ _3154_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__nor2_2
XFILLER_0_75_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5091_ _0497_ _0498_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__and2_4
X_4111_ _2620_ _1920_ _3131_ VGND VGND VPWR VPWR _3219_ sky130_fd_sc_hd__mux2_1
X_4042_ _3149_ _3150_ _0947_ VGND VGND VPWR VPWR _3151_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5993_ _1483_ _1484_ _0991_ net48 VGND VGND VPWR VPWR _1485_ sky130_fd_sc_hd__and4b_1
XFILLER_0_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4944_ net36 VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_19_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4875_ _0261_ _0262_ _0253_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6614_ _2151_ _2152_ _2162_ VGND VGND VPWR VPWR _2164_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_74_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3826_ _0357_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3757_ _0281_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6545_ _2056_ _2087_ _2088_ VGND VGND VPWR VPWR _2089_ sky130_fd_sc_hd__nand3_1
XFILLER_0_43_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6476_ _1874_ _1877_ VGND VGND VPWR VPWR _2013_ sky130_fd_sc_hd__or2_2
XFILLER_0_42_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5427_ _0429_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5358_ _0788_ _0789_ _0790_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__nand3_1
XFILLER_0_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4309_ _3414_ _3387_ _3388_ net123 _3162_ VGND VGND VPWR VPWR _3415_ sky130_fd_sc_hd__a221o_1
X_5289_ _0699_ _0700_ _0715_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__o21ba_2
X_7028_ _0357_ _1056_ net52 net53 VGND VGND VPWR VPWR _2617_ sky130_fd_sc_hd__and4_1
XFILLER_0_69_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_694 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4660_ _3624_ _0028_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6330_ _0390_ net17 net18 _0488_ VGND VGND VPWR VPWR _1853_ sky130_fd_sc_hd__a22o_1
X_4591_ _3573_ _3601_ _3688_ VGND VGND VPWR VPWR _3694_ sky130_fd_sc_hd__or3b_1
XFILLER_0_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6261_ _1299_ _1777_ _1446_ VGND VGND VPWR VPWR _1779_ sky130_fd_sc_hd__a21oi_1
X_6192_ net178 net16 net17 _3242_ VGND VGND VPWR VPWR _1703_ sky130_fd_sc_hd__a22o_1
X_5212_ _3451_ _3452_ _2489_ _2521_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__nand4_2
X_5143_ _0546_ _0555_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5074_ _0476_ _0478_ _0479_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4025_ _2762_ VGND VGND VPWR VPWR _3134_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5976_ _1963_ _1942_ _1909_ _1876_ _0863_ _0864_ VGND VGND VPWR VPWR _1466_ sky130_fd_sc_hd__mux4_1
XFILLER_0_118_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4927_ _3305_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4858_ _0239_ _0244_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_7_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3809_ _0838_ _0849_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__nand2_4
XFILLER_0_7_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4789_ _0168_ _0169_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6528_ _2061_ _2069_ VGND VGND VPWR VPWR _2070_ sky130_fd_sc_hd__xor2_2
X_6459_ _0303_ net17 VGND VGND VPWR VPWR _1994_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5830_ _1299_ _1305_ VGND VGND VPWR VPWR _1306_ sky130_fd_sc_hd__xnor2_1
X_5761_ _1229_ _1230_ VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__xor2_1
XFILLER_0_56_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4712_ _0084_ _0086_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7431_ _0455_ _0696_ VGND VGND VPWR VPWR _3057_ sky130_fd_sc_hd__nand2_1
X_5692_ _1063_ _1065_ VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4643_ _3688_ _3690_ _0011_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4574_ _3674_ _3675_ _3612_ VGND VGND VPWR VPWR _3677_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7362_ _0293_ _3128_ VGND VGND VPWR VPWR _2982_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7293_ _2902_ _2905_ VGND VGND VPWR VPWR _2906_ sky130_fd_sc_hd__xor2_1
X_6313_ _2117_ _0654_ _1831_ _1833_ VGND VGND VPWR VPWR _1835_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_12_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6244_ _0428_ _3410_ VGND VGND VPWR VPWR _1760_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6175_ _2215_ _0219_ _1682_ _1683_ VGND VGND VPWR VPWR _1684_ sky130_fd_sc_hd__nand4_2
X_5126_ _0447_ _0408_ _0536_ _0537_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__a211o_1
X_5057_ _0450_ _0460_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4008_ _3024_ VGND VGND VPWR VPWR _3035_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5959_ _1446_ VGND VGND VPWR VPWR _1447_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_4 _3228_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4290_ _3159_ _2991_ _3215_ _3276_ _2914_ VGND VGND VPWR VPWR _3396_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_67_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer27 net150 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_1
Xrebuffer16 _0679_ VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__buf_1
Xrebuffer49 _0396_ VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__dlygate4sd1_1
X_6931_ _2507_ _2508_ _2509_ VGND VGND VPWR VPWR _2511_ sky130_fd_sc_hd__nand3_1
XFILLER_0_88_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_815 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer38 _1255_ VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__dlygate4sd1_1
X_6862_ _2185_ _2187_ _2433_ _2435_ VGND VGND VPWR VPWR _2436_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5813_ _1021_ _1029_ _1272_ VGND VGND VPWR VPWR _1289_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6793_ _3386_ _1865_ _2358_ _2359_ VGND VGND VPWR VPWR _2360_ sky130_fd_sc_hd__nand4_1
XFILLER_0_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5744_ _1195_ _1196_ _1212_ VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__o21a_2
XFILLER_0_57_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5675_ net134 _1136_ _1137_ VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__nand3_2
XFILLER_0_60_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4626_ _1843_ _1985_ _2631_ _2806_ _3087_ _3301_ VGND VGND VPWR VPWR _3728_ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7414_ _3029_ _3038_ VGND VGND VPWR VPWR _3039_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7345_ _2961_ _2962_ VGND VGND VPWR VPWR _2963_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4557_ _3657_ _3658_ _3649_ VGND VGND VPWR VPWR _3660_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4488_ _3490_ _3591_ _3486_ VGND VGND VPWR VPWR _3592_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7276_ net56 _2051_ VGND VGND VPWR VPWR _2887_ sky130_fd_sc_hd__or2b_1
XFILLER_0_40_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6227_ _1678_ _1680_ _1739_ _1740_ VGND VGND VPWR VPWR _1741_ sky130_fd_sc_hd__or4_4
X_6158_ _2445_ _0688_ _1662_ _1663_ VGND VGND VPWR VPWR _1665_ sky130_fd_sc_hd__a22o_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _0516_ _0517_ _0518_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__nand3_4
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6089_ _1588_ _1589_ VGND VGND VPWR VPWR _1590_ sky130_fd_sc_hd__nand2_2
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput85 net167 VGND VGND VPWR VPWR result[24] sky130_fd_sc_hd__clkbuf_4
Xoutput74 net74 VGND VGND VPWR VPWR result[14] sky130_fd_sc_hd__clkbuf_4
Xoutput96 net96 VGND VGND VPWR VPWR result[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_829 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3790_ _0630_ _0641_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__nor2_4
XFILLER_0_109_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5460_ _0707_ _0466_ _0721_ _0874_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__and4_1
XFILLER_0_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4411_ _0707_ _0477_ _3424_ _3512_ VGND VGND VPWR VPWR _3515_ sky130_fd_sc_hd__and4_2
XFILLER_0_151_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5391_ _2587_ _0722_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4342_ _0292_ _2423_ VGND VGND VPWR VPWR _3447_ sky130_fd_sc_hd__and2_1
X_7130_ _2903_ _1745_ _2515_ _2514_ VGND VGND VPWR VPWR _2728_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4273_ _3257_ _3334_ _3377_ _3378_ VGND VGND VPWR VPWR _3379_ sky130_fd_sc_hd__or4_4
X_7061_ _2502_ _2481_ _2651_ _2652_ VGND VGND VPWR VPWR _2654_ sky130_fd_sc_hd__o211a_1
X_6012_ _2390_ _0654_ _1502_ _1503_ VGND VGND VPWR VPWR _1506_ sky130_fd_sc_hd__a22o_1
.ends


module alu_32_bit (zero_flag,
    A,
    B,
    control,
    result);
 output zero_flag;
 input [31:0] A;
 input [31:0] B;
 input [3:0] control;
 output [31:0] result;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;

 sky130_fd_sc_hd__buf_6 _3733_ (.A(net59),
    .X(_0030_));
 sky130_fd_sc_hd__buf_6 _3734_ (.A(_0030_),
    .X(_0041_));
 sky130_fd_sc_hd__buf_6 _3735_ (.A(_0041_),
    .X(_0052_));
 sky130_fd_sc_hd__clkbuf_4 _3736_ (.A(_0052_),
    .X(_0063_));
 sky130_fd_sc_hd__buf_6 _3737_ (.A(net27),
    .X(_0074_));
 sky130_fd_sc_hd__buf_2 _3738_ (.A(_0074_),
    .X(_0085_));
 sky130_fd_sc_hd__buf_4 _3739_ (.A(_0085_),
    .X(_0095_));
 sky130_fd_sc_hd__buf_6 _3740_ (.A(_0095_),
    .X(_0106_));
 sky130_fd_sc_hd__buf_6 _3741_ (.A(_0106_),
    .X(_0117_));
 sky130_fd_sc_hd__and2_1 _3742_ (.A(_0063_),
    .B(_0117_),
    .X(_0128_));
 sky130_fd_sc_hd__nor2_1 _3743_ (.A(_0063_),
    .B(_0117_),
    .Y(_0139_));
 sky130_fd_sc_hd__or2_1 _3744_ (.A(_0128_),
    .B(_0139_),
    .X(_0150_));
 sky130_fd_sc_hd__buf_6 _3745_ (.A(net58),
    .X(_0161_));
 sky130_fd_sc_hd__buf_4 _3746_ (.A(_0161_),
    .X(_0172_));
 sky130_fd_sc_hd__clkbuf_4 _3747_ (.A(_0172_),
    .X(_0183_));
 sky130_fd_sc_hd__clkbuf_4 _3748_ (.A(net26),
    .X(_0194_));
 sky130_fd_sc_hd__buf_4 _3749_ (.A(_0194_),
    .X(_0205_));
 sky130_fd_sc_hd__clkbuf_4 _3750_ (.A(_0205_),
    .X(_0215_));
 sky130_fd_sc_hd__buf_4 _3751_ (.A(_0215_),
    .X(_0226_));
 sky130_fd_sc_hd__nand2_1 _3752_ (.A(_0183_),
    .B(_0226_),
    .Y(_0237_));
 sky130_fd_sc_hd__or2_1 _3753_ (.A(_0183_),
    .B(_0226_),
    .X(_0248_));
 sky130_fd_sc_hd__nand2_1 _3754_ (.A(_0237_),
    .B(_0248_),
    .Y(_0259_));
 sky130_fd_sc_hd__and2_1 _3755_ (.A(net55),
    .B(net23),
    .X(_0270_));
 sky130_fd_sc_hd__buf_4 _3756_ (.A(net55),
    .X(_0281_));
 sky130_fd_sc_hd__buf_2 _3757_ (.A(_0281_),
    .X(_0292_));
 sky130_fd_sc_hd__buf_4 _3758_ (.A(_0292_),
    .X(_0303_));
 sky130_fd_sc_hd__buf_6 _3759_ (.A(net23),
    .X(_0314_));
 sky130_fd_sc_hd__buf_6 _3760_ (.A(_0314_),
    .X(_0324_));
 sky130_fd_sc_hd__clkbuf_4 _3761_ (.A(_0324_),
    .X(_0335_));
 sky130_fd_sc_hd__clkbuf_4 _3762_ (.A(_0335_),
    .X(_0346_));
 sky130_fd_sc_hd__buf_4 _3763_ (.A(_0346_),
    .X(_0357_));
 sky130_fd_sc_hd__nor2_1 _3764_ (.A(_0303_),
    .B(_0357_),
    .Y(_0368_));
 sky130_fd_sc_hd__or2_2 _3765_ (.A(_0270_),
    .B(_0368_),
    .X(_0379_));
 sky130_fd_sc_hd__clkbuf_4 _3766_ (.A(net44),
    .X(_0390_));
 sky130_fd_sc_hd__buf_4 _3767_ (.A(_0390_),
    .X(_0401_));
 sky130_fd_sc_hd__buf_6 _3768_ (.A(net12),
    .X(_0412_));
 sky130_fd_sc_hd__buf_2 _3769_ (.A(_0412_),
    .X(_0423_));
 sky130_fd_sc_hd__buf_4 _3770_ (.A(_0423_),
    .X(_0434_));
 sky130_fd_sc_hd__buf_4 _3771_ (.A(_0434_),
    .X(_0445_));
 sky130_fd_sc_hd__xnor2_2 _3772_ (.A(_0401_),
    .B(_0445_),
    .Y(_0455_));
 sky130_fd_sc_hd__clkbuf_4 _3773_ (.A(net1),
    .X(_0466_));
 sky130_fd_sc_hd__buf_4 _3774_ (.A(_0466_),
    .X(_0477_));
 sky130_fd_sc_hd__clkbuf_4 _3775_ (.A(net33),
    .X(_0488_));
 sky130_fd_sc_hd__buf_4 _3776_ (.A(_0488_),
    .X(_0499_));
 sky130_fd_sc_hd__or2b_2 _3777_ (.A(_0477_),
    .B_N(_0499_),
    .X(_0510_));
 sky130_fd_sc_hd__clkbuf_4 _3778_ (.A(_0401_),
    .X(_0521_));
 sky130_fd_sc_hd__and2b_1 _3779_ (.A_N(_0521_),
    .B(_0445_),
    .X(_0532_));
 sky130_fd_sc_hd__a21o_1 _3780_ (.A1(_0455_),
    .A2(_0510_),
    .B1(_0532_),
    .X(_0543_));
 sky130_fd_sc_hd__inv_2 _3781_ (.A(_0303_),
    .Y(_0554_));
 sky130_fd_sc_hd__and2_1 _3782_ (.A(_0554_),
    .B(_0357_),
    .X(_0565_));
 sky130_fd_sc_hd__a21o_1 _3783_ (.A1(_0379_),
    .A2(_0543_),
    .B1(_0565_),
    .X(_0576_));
 sky130_fd_sc_hd__inv_2 _3784_ (.A(_0172_),
    .Y(_0587_));
 sky130_fd_sc_hd__and2_1 _3785_ (.A(_0587_),
    .B(_0226_),
    .X(_0597_));
 sky130_fd_sc_hd__a21o_1 _3786_ (.A1(_0259_),
    .A2(_0576_),
    .B1(_0597_),
    .X(_0608_));
 sky130_fd_sc_hd__or2_1 _3787_ (.A(_0150_),
    .B(_0608_),
    .X(_0619_));
 sky130_fd_sc_hd__inv_2 _3788_ (.A(net65),
    .Y(_0630_));
 sky130_fd_sc_hd__or3_4 _3789_ (.A(net66),
    .B(net67),
    .C(net68),
    .X(_0641_));
 sky130_fd_sc_hd__nor2_4 _3790_ (.A(_0630_),
    .B(_0641_),
    .Y(_0652_));
 sky130_fd_sc_hd__nand2_1 _3791_ (.A(_0150_),
    .B(_0608_),
    .Y(_0663_));
 sky130_fd_sc_hd__nor2_1 _3792_ (.A(_0183_),
    .B(_0226_),
    .Y(_0674_));
 sky130_fd_sc_hd__nor2_1 _3793_ (.A(_0521_),
    .B(_0445_),
    .Y(_0685_));
 sky130_fd_sc_hd__nand2_2 _3794_ (.A(_0499_),
    .B(_0477_),
    .Y(_0696_));
 sky130_fd_sc_hd__buf_4 _3795_ (.A(_0423_),
    .X(_0707_));
 sky130_fd_sc_hd__and2_1 _3796_ (.A(_0401_),
    .B(_0707_),
    .X(_0717_));
 sky130_fd_sc_hd__o21ba_1 _3797_ (.A1(_0685_),
    .A2(_0696_),
    .B1_N(_0717_),
    .X(_0728_));
 sky130_fd_sc_hd__buf_6 _3798_ (.A(_0324_),
    .X(_0739_));
 sky130_fd_sc_hd__nand2_2 _3799_ (.A(_0303_),
    .B(_0739_),
    .Y(_0750_));
 sky130_fd_sc_hd__o21a_1 _3800_ (.A1(_0368_),
    .A2(_0728_),
    .B1(_0750_),
    .X(_0761_));
 sky130_fd_sc_hd__o21a_1 _3801_ (.A1(_0674_),
    .A2(_0761_),
    .B1(_0237_),
    .X(_0772_));
 sky130_fd_sc_hd__clkbuf_4 _3802_ (.A(net65),
    .X(_0783_));
 sky130_fd_sc_hd__nor2_1 _3803_ (.A(_0783_),
    .B(_0641_),
    .Y(_0794_));
 sky130_fd_sc_hd__o21ai_1 _3804_ (.A1(_0150_),
    .A2(_0772_),
    .B1(_0794_),
    .Y(_0805_));
 sky130_fd_sc_hd__a21oi_1 _3805_ (.A1(_0150_),
    .A2(_0772_),
    .B1(_0805_),
    .Y(_0816_));
 sky130_fd_sc_hd__inv_2 _3806_ (.A(_0052_),
    .Y(_0827_));
 sky130_fd_sc_hd__buf_4 _3807_ (.A(_0827_),
    .X(_0838_));
 sky130_fd_sc_hd__and4bb_4 _3808_ (.A_N(net66),
    .B_N(net68),
    .C(net67),
    .D(net65),
    .X(_0849_));
 sky130_fd_sc_hd__nand2_4 _3809_ (.A(_0838_),
    .B(_0849_),
    .Y(_0860_));
 sky130_fd_sc_hd__buf_2 _3810_ (.A(_0183_),
    .X(_0870_));
 sky130_fd_sc_hd__clkbuf_4 _3811_ (.A(_0499_),
    .X(_0881_));
 sky130_fd_sc_hd__buf_4 _3812_ (.A(_0881_),
    .X(_0892_));
 sky130_fd_sc_hd__clkbuf_4 _3813_ (.A(_0892_),
    .X(_0903_));
 sky130_fd_sc_hd__buf_4 _3814_ (.A(_0903_),
    .X(_0914_));
 sky130_fd_sc_hd__clkbuf_4 _3815_ (.A(_0914_),
    .X(_0925_));
 sky130_fd_sc_hd__clkbuf_4 _3816_ (.A(_0521_),
    .X(_0936_));
 sky130_fd_sc_hd__clkbuf_4 _3817_ (.A(_0936_),
    .X(_0947_));
 sky130_fd_sc_hd__clkbuf_4 _3818_ (.A(_0947_),
    .X(_0958_));
 sky130_fd_sc_hd__clkbuf_4 _3819_ (.A(_0958_),
    .X(_0969_));
 sky130_fd_sc_hd__clkbuf_4 _3820_ (.A(_0303_),
    .X(_0980_));
 sky130_fd_sc_hd__clkbuf_4 _3821_ (.A(_0466_),
    .X(_0991_));
 sky130_fd_sc_hd__buf_4 _3822_ (.A(_0991_),
    .X(_1002_));
 sky130_fd_sc_hd__nand2_2 _3823_ (.A(_0980_),
    .B(_1002_),
    .Y(_1012_));
 sky130_fd_sc_hd__buf_4 _3824_ (.A(_0117_),
    .X(_1023_));
 sky130_fd_sc_hd__buf_4 _3825_ (.A(_0226_),
    .X(_1034_));
 sky130_fd_sc_hd__clkbuf_4 _3826_ (.A(_0357_),
    .X(_1045_));
 sky130_fd_sc_hd__buf_4 _3827_ (.A(_0445_),
    .X(_1056_));
 sky130_fd_sc_hd__buf_4 _3828_ (.A(_1056_),
    .X(_1067_));
 sky130_fd_sc_hd__mux4_1 _3829_ (.A0(_1023_),
    .A1(_1034_),
    .A2(_1045_),
    .A3(_1067_),
    .S0(_0903_),
    .S1(_0947_),
    .X(_1078_));
 sky130_fd_sc_hd__inv_2 _3830_ (.A(_1078_),
    .Y(_1089_));
 sky130_fd_sc_hd__clkbuf_4 _3831_ (.A(_0980_),
    .X(_1100_));
 sky130_fd_sc_hd__o32a_1 _3832_ (.A1(_0925_),
    .A2(_0969_),
    .A3(_1012_),
    .B1(_1089_),
    .B2(_1100_),
    .X(_1111_));
 sky130_fd_sc_hd__or2_1 _3833_ (.A(_0870_),
    .B(_1111_),
    .X(_1122_));
 sky130_fd_sc_hd__nor2_1 _3834_ (.A(_0860_),
    .B(_1122_),
    .Y(_1133_));
 sky130_fd_sc_hd__buf_2 _3835_ (.A(net67),
    .X(_1144_));
 sky130_fd_sc_hd__clkbuf_2 _3836_ (.A(net68),
    .X(_1154_));
 sky130_fd_sc_hd__clkbuf_2 _3837_ (.A(net66),
    .X(_1165_));
 sky130_fd_sc_hd__nor4b_2 _3838_ (.A(_0783_),
    .B(_1144_),
    .C(_1154_),
    .D_N(_1165_),
    .Y(_1176_));
 sky130_fd_sc_hd__and4bb_2 _3839_ (.A_N(_1165_),
    .B_N(_1144_),
    .C(_1154_),
    .D(net65),
    .X(_1187_));
 sky130_fd_sc_hd__or4b_1 _3840_ (.A(net66),
    .B(net65),
    .C(net68),
    .D_N(net67),
    .X(_1198_));
 sky130_fd_sc_hd__buf_2 _3841_ (.A(_1198_),
    .X(_1209_));
 sky130_fd_sc_hd__and4bb_2 _3842_ (.A_N(_1144_),
    .B_N(_1154_),
    .C(_1165_),
    .D(net65),
    .X(_1220_));
 sky130_fd_sc_hd__o21ba_1 _3843_ (.A1(_0128_),
    .A2(_1209_),
    .B1_N(_1220_),
    .X(_1231_));
 sky130_fd_sc_hd__nor2_1 _3844_ (.A(_0139_),
    .B(_1231_),
    .Y(_1242_));
 sky130_fd_sc_hd__a221o_1 _3845_ (.A1(_0128_),
    .A2(_1176_),
    .B1(_1187_),
    .B2(_0139_),
    .C1(_1242_),
    .X(_1253_));
 sky130_fd_sc_hd__clkbuf_4 _3846_ (.A(net26),
    .X(_1264_));
 sky130_fd_sc_hd__clkbuf_4 _3847_ (.A(_1264_),
    .X(_1275_));
 sky130_fd_sc_hd__and4_1 _3848_ (.A(_1275_),
    .B(_0499_),
    .C(_0401_),
    .D(_0739_),
    .X(_1286_));
 sky130_fd_sc_hd__a22o_1 _3849_ (.A1(_1275_),
    .A2(_0499_),
    .B1(_0401_),
    .B2(_0739_),
    .X(_1296_));
 sky130_fd_sc_hd__or2b_1 _3850_ (.A(_1286_),
    .B_N(_1296_),
    .X(_1307_));
 sky130_fd_sc_hd__nand2_1 _3851_ (.A(_0303_),
    .B(_0445_),
    .Y(_1318_));
 sky130_fd_sc_hd__xnor2_1 _3852_ (.A(_1307_),
    .B(_1318_),
    .Y(_1329_));
 sky130_fd_sc_hd__a21o_1 _3853_ (.A1(_0881_),
    .A2(_0357_),
    .B1(_0717_),
    .X(_1340_));
 sky130_fd_sc_hd__and3_1 _3854_ (.A(_0881_),
    .B(_0357_),
    .C(_0717_),
    .X(_1351_));
 sky130_fd_sc_hd__a31o_1 _3855_ (.A1(_0980_),
    .A2(_1002_),
    .A3(_1340_),
    .B1(_1351_),
    .X(_1362_));
 sky130_fd_sc_hd__or2b_1 _3856_ (.A(_1329_),
    .B_N(_1362_),
    .X(_1373_));
 sky130_fd_sc_hd__buf_4 _3857_ (.A(_1002_),
    .X(_1384_));
 sky130_fd_sc_hd__xnor2_1 _3858_ (.A(_1329_),
    .B(_1362_),
    .Y(_1395_));
 sky130_fd_sc_hd__nand3_1 _3859_ (.A(_0183_),
    .B(_1384_),
    .C(_1395_),
    .Y(_1406_));
 sky130_fd_sc_hd__a22o_1 _3860_ (.A1(_0172_),
    .A2(_0707_),
    .B1(_0477_),
    .B2(_0052_),
    .X(_1417_));
 sky130_fd_sc_hd__inv_2 _3861_ (.A(_0423_),
    .Y(_1428_));
 sky130_fd_sc_hd__or4b_4 _3862_ (.A(_0587_),
    .B(_0827_),
    .C(_1428_),
    .D_N(_0466_),
    .X(_1439_));
 sky130_fd_sc_hd__a31o_1 _3863_ (.A1(_0303_),
    .A2(_0434_),
    .A3(_1296_),
    .B1(_1286_),
    .X(_1449_));
 sky130_fd_sc_hd__and4_1 _3864_ (.A(net194),
    .B(net26),
    .C(net33),
    .D(net44),
    .X(_1460_));
 sky130_fd_sc_hd__a22o_1 _3865_ (.A1(net194),
    .A2(net33),
    .B1(net44),
    .B2(net26),
    .X(_1471_));
 sky130_fd_sc_hd__and2b_1 _3866_ (.A_N(_1460_),
    .B(_1471_),
    .X(_1482_));
 sky130_fd_sc_hd__xnor2_1 _3867_ (.A(_0750_),
    .B(_1482_),
    .Y(_1493_));
 sky130_fd_sc_hd__xor2_1 _3868_ (.A(_1449_),
    .B(_1493_),
    .X(_1504_));
 sky130_fd_sc_hd__and3_1 _3869_ (.A(_1417_),
    .B(_1439_),
    .C(_1504_),
    .X(_1515_));
 sky130_fd_sc_hd__a21oi_1 _3870_ (.A1(_1417_),
    .A2(_1439_),
    .B1(_1504_),
    .Y(_1526_));
 sky130_fd_sc_hd__or2_1 _3871_ (.A(_1515_),
    .B(_1526_),
    .X(_1537_));
 sky130_fd_sc_hd__a21o_1 _3872_ (.A1(_1373_),
    .A2(_1406_),
    .B1(_1537_),
    .X(_1548_));
 sky130_fd_sc_hd__nand3_1 _3873_ (.A(_1373_),
    .B(_1406_),
    .C(_1537_),
    .Y(_1559_));
 sky130_fd_sc_hd__and2_1 _3874_ (.A(_1548_),
    .B(_1559_),
    .X(_1570_));
 sky130_fd_sc_hd__and2b_1 _3875_ (.A_N(_1351_),
    .B(_1340_),
    .X(_1581_));
 sky130_fd_sc_hd__xnor2_1 _3876_ (.A(_1012_),
    .B(_1581_),
    .Y(_1592_));
 sky130_fd_sc_hd__and4_1 _3877_ (.A(_0881_),
    .B(_0521_),
    .C(_1056_),
    .D(_1002_),
    .X(_1603_));
 sky130_fd_sc_hd__and2_1 _3878_ (.A(_1592_),
    .B(_1603_),
    .X(_1613_));
 sky130_fd_sc_hd__a21o_1 _3879_ (.A1(_0183_),
    .A2(_1384_),
    .B1(_1395_),
    .X(_1624_));
 sky130_fd_sc_hd__and2_1 _3880_ (.A(_1406_),
    .B(_1624_),
    .X(_1635_));
 sky130_fd_sc_hd__and2_1 _3881_ (.A(_1613_),
    .B(_1635_),
    .X(_1646_));
 sky130_fd_sc_hd__nand2_1 _3882_ (.A(_1570_),
    .B(_1646_),
    .Y(_1657_));
 sky130_fd_sc_hd__and4bb_2 _3883_ (.A_N(_0783_),
    .B_N(_1144_),
    .C(_1154_),
    .D(_1165_),
    .X(_1668_));
 sky130_fd_sc_hd__or2_1 _3884_ (.A(_1570_),
    .B(_1646_),
    .X(_1679_));
 sky130_fd_sc_hd__and3b_1 _3885_ (.A_N(net68),
    .B(net67),
    .C(net66),
    .X(_1690_));
 sky130_fd_sc_hd__buf_2 _3886_ (.A(_1690_),
    .X(_1701_));
 sky130_fd_sc_hd__clkbuf_4 _3887_ (.A(_0554_),
    .X(_1712_));
 sky130_fd_sc_hd__clkbuf_4 _3888_ (.A(_0587_),
    .X(_1723_));
 sky130_fd_sc_hd__nor2_2 _3889_ (.A(_1712_),
    .B(_1723_),
    .Y(_1734_));
 sky130_fd_sc_hd__buf_2 _3890_ (.A(net17),
    .X(_1745_));
 sky130_fd_sc_hd__buf_4 _3891_ (.A(_1745_),
    .X(_1756_));
 sky130_fd_sc_hd__buf_2 _3892_ (.A(net18),
    .X(_1767_));
 sky130_fd_sc_hd__buf_4 _3893_ (.A(_1767_),
    .X(_1778_));
 sky130_fd_sc_hd__mux2_1 _3894_ (.A0(_1756_),
    .A1(_1778_),
    .S(_0892_),
    .X(_1788_));
 sky130_fd_sc_hd__buf_2 _3895_ (.A(net19),
    .X(_1799_));
 sky130_fd_sc_hd__clkbuf_4 _3896_ (.A(_1799_),
    .X(_1810_));
 sky130_fd_sc_hd__clkbuf_4 _3897_ (.A(net20),
    .X(_1821_));
 sky130_fd_sc_hd__mux2_1 _3898_ (.A0(_1810_),
    .A1(_1821_),
    .S(_0892_),
    .X(_1832_));
 sky130_fd_sc_hd__mux2_1 _3899_ (.A0(_1788_),
    .A1(_1832_),
    .S(_0936_),
    .X(_1843_));
 sky130_fd_sc_hd__clkbuf_4 _3900_ (.A(net13),
    .X(_1854_));
 sky130_fd_sc_hd__buf_4 _3901_ (.A(_1854_),
    .X(_1865_));
 sky130_fd_sc_hd__clkbuf_4 _3902_ (.A(_1865_),
    .X(_1876_));
 sky130_fd_sc_hd__clkbuf_4 _3903_ (.A(net14),
    .X(_1887_));
 sky130_fd_sc_hd__clkbuf_4 _3904_ (.A(_1887_),
    .X(_1898_));
 sky130_fd_sc_hd__buf_4 _3905_ (.A(_1898_),
    .X(_1909_));
 sky130_fd_sc_hd__mux2_1 _3906_ (.A0(_1876_),
    .A1(_1909_),
    .S(_0892_),
    .X(_1920_));
 sky130_fd_sc_hd__clkbuf_4 _3907_ (.A(net15),
    .X(_1931_));
 sky130_fd_sc_hd__clkbuf_4 _3908_ (.A(_1931_),
    .X(_1942_));
 sky130_fd_sc_hd__buf_2 _3909_ (.A(net16),
    .X(_1952_));
 sky130_fd_sc_hd__buf_4 _3910_ (.A(_1952_),
    .X(_1963_));
 sky130_fd_sc_hd__mux2_1 _3911_ (.A0(_1942_),
    .A1(_1963_),
    .S(_0892_),
    .X(_1974_));
 sky130_fd_sc_hd__mux2_1 _3912_ (.A0(_1920_),
    .A1(_1974_),
    .S(_0936_),
    .X(_1985_));
 sky130_fd_sc_hd__mux2_1 _3913_ (.A0(_1843_),
    .A1(_1985_),
    .S(_0554_),
    .X(_1996_));
 sky130_fd_sc_hd__clkbuf_4 _3914_ (.A(net21),
    .X(_2007_));
 sky130_fd_sc_hd__clkbuf_4 _3915_ (.A(net22),
    .X(_2018_));
 sky130_fd_sc_hd__buf_6 _3916_ (.A(_0881_),
    .X(_2029_));
 sky130_fd_sc_hd__mux2_1 _3917_ (.A0(_2007_),
    .A1(_2018_),
    .S(_2029_),
    .X(_2040_));
 sky130_fd_sc_hd__clkbuf_4 _3918_ (.A(net24),
    .X(_2051_));
 sky130_fd_sc_hd__mux2_2 _3919_ (.A0(_2051_),
    .A1(net25),
    .S(_0892_),
    .X(_2062_));
 sky130_fd_sc_hd__mux2_2 _3920_ (.A0(_2040_),
    .A1(_2062_),
    .S(_0936_),
    .X(_2073_));
 sky130_fd_sc_hd__a21o_1 _3921_ (.A1(_0554_),
    .A2(_2073_),
    .B1(_0587_),
    .X(_2084_));
 sky130_fd_sc_hd__o21a_2 _3922_ (.A1(_0870_),
    .A2(_1996_),
    .B1(_2084_),
    .X(_2095_));
 sky130_fd_sc_hd__buf_4 _3923_ (.A(net31),
    .X(_2106_));
 sky130_fd_sc_hd__clkbuf_4 _3924_ (.A(_2106_),
    .X(_2117_));
 sky130_fd_sc_hd__clkbuf_4 _3925_ (.A(_2117_),
    .X(_2127_));
 sky130_fd_sc_hd__clkbuf_4 _3926_ (.A(_2127_),
    .X(_2138_));
 sky130_fd_sc_hd__buf_4 _3927_ (.A(net32),
    .X(_2149_));
 sky130_fd_sc_hd__clkbuf_4 _3928_ (.A(_2149_),
    .X(_2160_));
 sky130_fd_sc_hd__clkbuf_4 _3929_ (.A(_2160_),
    .X(_2171_));
 sky130_fd_sc_hd__clkbuf_4 _3930_ (.A(_2171_),
    .X(_2182_));
 sky130_fd_sc_hd__mux2_1 _3931_ (.A0(_2138_),
    .A1(_2182_),
    .S(_2029_),
    .X(_2193_));
 sky130_fd_sc_hd__clkbuf_4 _3932_ (.A(net2),
    .X(_2204_));
 sky130_fd_sc_hd__clkbuf_4 _3933_ (.A(_2204_),
    .X(_2215_));
 sky130_fd_sc_hd__buf_2 _3934_ (.A(_2215_),
    .X(_2226_));
 sky130_fd_sc_hd__clkbuf_4 _3935_ (.A(_2226_),
    .X(_2237_));
 sky130_fd_sc_hd__clkbuf_4 _3936_ (.A(net3),
    .X(_2248_));
 sky130_fd_sc_hd__clkbuf_4 _3937_ (.A(_2248_),
    .X(_2259_));
 sky130_fd_sc_hd__buf_4 _3938_ (.A(_2259_),
    .X(_2270_));
 sky130_fd_sc_hd__mux2_1 _3939_ (.A0(_2237_),
    .A1(_2270_),
    .S(_2029_),
    .X(_2281_));
 sky130_fd_sc_hd__mux2_1 _3940_ (.A0(_2193_),
    .A1(_2281_),
    .S(_0936_),
    .X(_2292_));
 sky130_fd_sc_hd__buf_4 _3941_ (.A(net28),
    .X(_2302_));
 sky130_fd_sc_hd__clkbuf_4 _3942_ (.A(_2302_),
    .X(_2313_));
 sky130_fd_sc_hd__buf_4 _3943_ (.A(_2313_),
    .X(_2324_));
 sky130_fd_sc_hd__buf_4 _3944_ (.A(_2324_),
    .X(_2335_));
 sky130_fd_sc_hd__buf_6 _3945_ (.A(_2335_),
    .X(_2346_));
 sky130_fd_sc_hd__mux2_1 _3946_ (.A0(_1023_),
    .A1(_2346_),
    .S(_2029_),
    .X(_2357_));
 sky130_fd_sc_hd__buf_4 _3947_ (.A(net29),
    .X(_2368_));
 sky130_fd_sc_hd__clkbuf_4 _3948_ (.A(_2368_),
    .X(_2379_));
 sky130_fd_sc_hd__buf_6 _3949_ (.A(_2379_),
    .X(_2390_));
 sky130_fd_sc_hd__buf_4 _3950_ (.A(_2390_),
    .X(_2401_));
 sky130_fd_sc_hd__buf_4 _3951_ (.A(_2401_),
    .X(_2412_));
 sky130_fd_sc_hd__buf_4 _3952_ (.A(net30),
    .X(_2423_));
 sky130_fd_sc_hd__buf_4 _3953_ (.A(_2423_),
    .X(_2434_));
 sky130_fd_sc_hd__buf_4 _3954_ (.A(_2434_),
    .X(_2445_));
 sky130_fd_sc_hd__clkbuf_4 _3955_ (.A(_2445_),
    .X(_2456_));
 sky130_fd_sc_hd__mux2_2 _3956_ (.A0(_2412_),
    .A1(_2456_),
    .S(_2029_),
    .X(_2467_));
 sky130_fd_sc_hd__mux2_1 _3957_ (.A0(_2357_),
    .A1(_2467_),
    .S(_0936_),
    .X(_2478_));
 sky130_fd_sc_hd__clkbuf_4 _3958_ (.A(net8),
    .X(_2489_));
 sky130_fd_sc_hd__clkbuf_4 _3959_ (.A(_2489_),
    .X(_2499_));
 sky130_fd_sc_hd__clkbuf_4 _3960_ (.A(_2499_),
    .X(_2510_));
 sky130_fd_sc_hd__clkbuf_4 _3961_ (.A(net9),
    .X(_2521_));
 sky130_fd_sc_hd__clkbuf_4 _3962_ (.A(_2521_),
    .X(_2532_));
 sky130_fd_sc_hd__clkbuf_4 _3963_ (.A(_2532_),
    .X(_2543_));
 sky130_fd_sc_hd__mux2_1 _3964_ (.A0(_2510_),
    .A1(_2543_),
    .S(_2029_),
    .X(_2554_));
 sky130_fd_sc_hd__buf_4 _3965_ (.A(net10),
    .X(_2565_));
 sky130_fd_sc_hd__clkbuf_4 _3966_ (.A(_2565_),
    .X(_2576_));
 sky130_fd_sc_hd__clkbuf_4 _3967_ (.A(_2576_),
    .X(_2587_));
 sky130_fd_sc_hd__clkbuf_4 _3968_ (.A(net11),
    .X(_2598_));
 sky130_fd_sc_hd__buf_4 _3969_ (.A(_2598_),
    .X(_2609_));
 sky130_fd_sc_hd__mux2_1 _3970_ (.A0(_2587_),
    .A1(_2609_),
    .S(_2029_),
    .X(_2620_));
 sky130_fd_sc_hd__mux2_1 _3971_ (.A0(_2554_),
    .A1(_2620_),
    .S(_0936_),
    .X(_2631_));
 sky130_fd_sc_hd__buf_4 _3972_ (.A(net4),
    .X(_2642_));
 sky130_fd_sc_hd__buf_4 _3973_ (.A(_2642_),
    .X(_2653_));
 sky130_fd_sc_hd__buf_4 _3974_ (.A(_2653_),
    .X(_2664_));
 sky130_fd_sc_hd__clkbuf_4 _3975_ (.A(_2664_),
    .X(_2675_));
 sky130_fd_sc_hd__buf_4 _3976_ (.A(net5),
    .X(_2686_));
 sky130_fd_sc_hd__buf_4 _3977_ (.A(_2686_),
    .X(_2696_));
 sky130_fd_sc_hd__buf_4 _3978_ (.A(_2696_),
    .X(_2707_));
 sky130_fd_sc_hd__buf_4 _3979_ (.A(_2707_),
    .X(_2718_));
 sky130_fd_sc_hd__mux2_1 _3980_ (.A0(_2675_),
    .A1(_2718_),
    .S(_2029_),
    .X(_2729_));
 sky130_fd_sc_hd__buf_4 _3981_ (.A(net6),
    .X(_2740_));
 sky130_fd_sc_hd__buf_4 _3982_ (.A(_2740_),
    .X(_2751_));
 sky130_fd_sc_hd__buf_4 _3983_ (.A(_2751_),
    .X(_2762_));
 sky130_fd_sc_hd__clkbuf_4 _3984_ (.A(net7),
    .X(_2773_));
 sky130_fd_sc_hd__buf_4 _3985_ (.A(_2773_),
    .X(_2784_));
 sky130_fd_sc_hd__mux2_1 _3986_ (.A0(_2762_),
    .A1(_2784_),
    .S(_2029_),
    .X(_2795_));
 sky130_fd_sc_hd__mux2_1 _3987_ (.A0(_2729_),
    .A1(_2795_),
    .S(_0936_),
    .X(_2806_));
 sky130_fd_sc_hd__mux4_1 _3988_ (.A0(_2292_),
    .A1(_2478_),
    .A2(_2631_),
    .A3(_2806_),
    .S0(_0554_),
    .S1(_0183_),
    .X(_2817_));
 sky130_fd_sc_hd__mux2_1 _3989_ (.A0(_2095_),
    .A1(_2817_),
    .S(_0838_),
    .X(_2828_));
 sky130_fd_sc_hd__a41o_1 _3990_ (.A1(_0063_),
    .A2(net25),
    .A3(_0783_),
    .A4(_1734_),
    .B1(_2828_),
    .X(_2839_));
 sky130_fd_sc_hd__a32o_1 _3991_ (.A1(_1657_),
    .A2(_1668_),
    .A3(_1679_),
    .B1(_1701_),
    .B2(_2839_),
    .X(_2850_));
 sky130_fd_sc_hd__or4_1 _3992_ (.A(_0816_),
    .B(_1133_),
    .C(_1253_),
    .D(_2850_),
    .X(_2861_));
 sky130_fd_sc_hd__a31o_1 _3993_ (.A1(_0619_),
    .A2(_0652_),
    .A3(_0663_),
    .B1(_2861_),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_4 _3994_ (.A(net60),
    .X(_2881_));
 sky130_fd_sc_hd__clkbuf_4 _3995_ (.A(_2881_),
    .X(_2892_));
 sky130_fd_sc_hd__clkbuf_4 _3996_ (.A(_2892_),
    .X(_2903_));
 sky130_fd_sc_hd__nor2_1 _3997_ (.A(_2335_),
    .B(_2903_),
    .Y(_2914_));
 sky130_fd_sc_hd__and2_2 _3998_ (.A(_2302_),
    .B(net60),
    .X(_2925_));
 sky130_fd_sc_hd__or2_1 _3999_ (.A(_2914_),
    .B(_2925_),
    .X(_2936_));
 sky130_fd_sc_hd__and2_1 _4000_ (.A(_0838_),
    .B(_0117_),
    .X(_2947_));
 sky130_fd_sc_hd__a21o_1 _4001_ (.A1(_0150_),
    .A2(_0608_),
    .B1(_2947_),
    .X(_2958_));
 sky130_fd_sc_hd__xor2_1 _4002_ (.A(_2936_),
    .B(_2958_),
    .X(_2969_));
 sky130_fd_sc_hd__clkbuf_4 _4003_ (.A(_0794_),
    .X(_2980_));
 sky130_fd_sc_hd__o21ba_1 _4004_ (.A1(_0139_),
    .A2(_0772_),
    .B1_N(_0128_),
    .X(_2991_));
 sky130_fd_sc_hd__or2_1 _4005_ (.A(_2936_),
    .B(_2991_),
    .X(_3002_));
 sky130_fd_sc_hd__nand2_1 _4006_ (.A(_2936_),
    .B(_2991_),
    .Y(_3013_));
 sky130_fd_sc_hd__nor2_1 _4007_ (.A(_0554_),
    .B(_0936_),
    .Y(_3024_));
 sky130_fd_sc_hd__inv_2 _4008_ (.A(_3024_),
    .Y(_3035_));
 sky130_fd_sc_hd__buf_4 _4009_ (.A(_0925_),
    .X(_3046_));
 sky130_fd_sc_hd__o21a_1 _4010_ (.A1(_3046_),
    .A2(_1428_),
    .B1(_0696_),
    .X(_3056_));
 sky130_fd_sc_hd__mux4_1 _4011_ (.A0(_2346_),
    .A1(_1034_),
    .A2(_1023_),
    .A3(_1045_),
    .S0(_0958_),
    .S1(_0925_),
    .X(_3066_));
 sky130_fd_sc_hd__clkbuf_4 _4012_ (.A(_1712_),
    .X(_3077_));
 sky130_fd_sc_hd__clkbuf_4 _4013_ (.A(_3077_),
    .X(_3087_));
 sky130_fd_sc_hd__a2bb2o_2 _4014_ (.A1_N(_3035_),
    .A2_N(_3056_),
    .B1(_3066_),
    .B2(_3087_),
    .X(_3097_));
 sky130_fd_sc_hd__buf_2 _4015_ (.A(_0870_),
    .X(_3108_));
 sky130_fd_sc_hd__or4b_4 _4016_ (.A(_1165_),
    .B(_0630_),
    .C(_1154_),
    .D_N(_1144_),
    .X(_3118_));
 sky130_fd_sc_hd__nor2_2 _4017_ (.A(_3108_),
    .B(_3118_),
    .Y(_3126_));
 sky130_fd_sc_hd__buf_2 _4018_ (.A(_0063_),
    .X(_3127_));
 sky130_fd_sc_hd__clkbuf_4 _4019_ (.A(_2543_),
    .X(_3128_));
 sky130_fd_sc_hd__mux2_1 _4020_ (.A0(_3128_),
    .A1(_2587_),
    .S(_0903_),
    .X(_3129_));
 sky130_fd_sc_hd__mux2_1 _4021_ (.A0(_2609_),
    .A1(_1865_),
    .S(_0892_),
    .X(_3130_));
 sky130_fd_sc_hd__buf_4 _4022_ (.A(_0947_),
    .X(_3131_));
 sky130_fd_sc_hd__mux2_1 _4023_ (.A0(_3129_),
    .A1(_3130_),
    .S(_3131_),
    .X(_3132_));
 sky130_fd_sc_hd__clkbuf_4 _4024_ (.A(_2718_),
    .X(_3133_));
 sky130_fd_sc_hd__clkbuf_4 _4025_ (.A(_2762_),
    .X(_3134_));
 sky130_fd_sc_hd__clkbuf_4 _4026_ (.A(_2784_),
    .X(_3135_));
 sky130_fd_sc_hd__mux4_2 _4027_ (.A0(_3133_),
    .A1(_3134_),
    .A2(_3135_),
    .A3(_2510_),
    .S0(_0914_),
    .S1(_0958_),
    .X(_3136_));
 sky130_fd_sc_hd__clkbuf_4 _4028_ (.A(_2270_),
    .X(_3137_));
 sky130_fd_sc_hd__mux4_1 _4029_ (.A0(_2182_),
    .A1(_2237_),
    .A2(_3137_),
    .A3(_2675_),
    .S0(_0914_),
    .S1(_0958_),
    .X(_3138_));
 sky130_fd_sc_hd__buf_4 _4030_ (.A(_2456_),
    .X(_3139_));
 sky130_fd_sc_hd__mux4_1 _4031_ (.A0(_2346_),
    .A1(_2412_),
    .A2(_3139_),
    .A3(_2138_),
    .S0(_0914_),
    .S1(_0958_),
    .X(_3140_));
 sky130_fd_sc_hd__mux4_1 _4032_ (.A0(_3132_),
    .A1(_3136_),
    .A2(_3138_),
    .A3(_3140_),
    .S0(_3077_),
    .S1(_1723_),
    .X(_3141_));
 sky130_fd_sc_hd__and2b_1 _4033_ (.A_N(_0903_),
    .B(_2018_),
    .X(_3142_));
 sky130_fd_sc_hd__a21oi_1 _4034_ (.A1(_0903_),
    .A2(_2051_),
    .B1(_3142_),
    .Y(_3143_));
 sky130_fd_sc_hd__or2b_2 _4035_ (.A(_0903_),
    .B_N(net25),
    .X(_3144_));
 sky130_fd_sc_hd__mux2_1 _4036_ (.A0(_3143_),
    .A1(_3144_),
    .S(_3131_),
    .X(_3145_));
 sky130_fd_sc_hd__mux2_1 _4037_ (.A0(_1767_),
    .A1(_1799_),
    .S(_0892_),
    .X(_3146_));
 sky130_fd_sc_hd__mux2_1 _4038_ (.A0(_1821_),
    .A1(_2007_),
    .S(_2029_),
    .X(_3147_));
 sky130_fd_sc_hd__mux2_1 _4039_ (.A0(_3146_),
    .A1(_3147_),
    .S(_0947_),
    .X(_3148_));
 sky130_fd_sc_hd__mux2_1 _4040_ (.A0(_1909_),
    .A1(_1942_),
    .S(_0892_),
    .X(_3149_));
 sky130_fd_sc_hd__mux2_1 _4041_ (.A0(_1952_),
    .A1(_1745_),
    .S(_0892_),
    .X(_3150_));
 sky130_fd_sc_hd__mux2_1 _4042_ (.A0(_3149_),
    .A1(_3150_),
    .S(_0947_),
    .X(_3151_));
 sky130_fd_sc_hd__mux2_1 _4043_ (.A0(_3148_),
    .A1(_3151_),
    .S(_1712_),
    .X(_3152_));
 sky130_fd_sc_hd__nor2_1 _4044_ (.A(_0870_),
    .B(_3152_),
    .Y(_3153_));
 sky130_fd_sc_hd__nand3b_2 _4045_ (.A_N(_1154_),
    .B(_1144_),
    .C(_1165_),
    .Y(_3154_));
 sky130_fd_sc_hd__a2111o_1 _4046_ (.A1(_3108_),
    .A2(_3145_),
    .B1(_3153_),
    .C1(_1734_),
    .D1(_3154_),
    .X(_3155_));
 sky130_fd_sc_hd__nand2_4 _4047_ (.A(_0838_),
    .B(_1701_),
    .Y(_3156_));
 sky130_fd_sc_hd__a2bb2oi_1 _4048_ (.A1_N(_3127_),
    .A2_N(_3141_),
    .B1(_3155_),
    .B2(_3156_),
    .Y(_3157_));
 sky130_fd_sc_hd__nor4b_2 _4049_ (.A(net66),
    .B(net65),
    .C(net68),
    .D_N(net67),
    .Y(_3158_));
 sky130_fd_sc_hd__nand2_1 _4050_ (.A(_2346_),
    .B(_2903_),
    .Y(_3159_));
 sky130_fd_sc_hd__a21oi_1 _4051_ (.A1(_3158_),
    .A2(_3159_),
    .B1(_1220_),
    .Y(_3160_));
 sky130_fd_sc_hd__and3_4 _4052_ (.A(net25),
    .B(net65),
    .C(_1701_),
    .X(_3161_));
 sky130_fd_sc_hd__and3_2 _4053_ (.A(_0870_),
    .B(_0063_),
    .C(_3161_),
    .X(_3162_));
 sky130_fd_sc_hd__a21o_1 _4054_ (.A1(_0925_),
    .A2(_0969_),
    .B1(_1100_),
    .X(_3163_));
 sky130_fd_sc_hd__a2bb2o_1 _4055_ (.A1_N(_2914_),
    .A2_N(_3160_),
    .B1(_3162_),
    .B2(_3163_),
    .X(_3164_));
 sky130_fd_sc_hd__a221o_1 _4056_ (.A1(_1187_),
    .A2(_2914_),
    .B1(_2925_),
    .B2(_1176_),
    .C1(_3164_),
    .X(_3165_));
 sky130_fd_sc_hd__a311o_1 _4057_ (.A1(_0838_),
    .A2(_3097_),
    .A3(_3126_),
    .B1(_3157_),
    .C1(_3165_),
    .X(_3166_));
 sky130_fd_sc_hd__a31o_1 _4058_ (.A1(_2980_),
    .A2(_3002_),
    .A3(_3013_),
    .B1(_3166_),
    .X(_3167_));
 sky130_fd_sc_hd__and2_1 _4059_ (.A(_1449_),
    .B(_1493_),
    .X(_3168_));
 sky130_fd_sc_hd__buf_4 _4060_ (.A(net58),
    .X(_3169_));
 sky130_fd_sc_hd__a22oi_1 _4061_ (.A1(_3169_),
    .A2(_0314_),
    .B1(_0412_),
    .B2(net191),
    .Y(_3170_));
 sky130_fd_sc_hd__and4_1 _4062_ (.A(net58),
    .B(net59),
    .C(net23),
    .D(net12),
    .X(_3171_));
 sky130_fd_sc_hd__nor2_1 _4063_ (.A(_3170_),
    .B(_3171_),
    .Y(_3172_));
 sky130_fd_sc_hd__nand2_1 _4064_ (.A(net1),
    .B(net60),
    .Y(_3173_));
 sky130_fd_sc_hd__xor2_2 _4065_ (.A(_3172_),
    .B(_3173_),
    .X(_3174_));
 sky130_fd_sc_hd__and2_1 _4066_ (.A(_0281_),
    .B(net26),
    .X(_3175_));
 sky130_fd_sc_hd__buf_6 _4067_ (.A(net44),
    .X(_3176_));
 sky130_fd_sc_hd__nand4_2 _4068_ (.A(net194),
    .B(net33),
    .C(_3176_),
    .D(net28),
    .Y(_3177_));
 sky130_fd_sc_hd__a22o_1 _4069_ (.A1(net194),
    .A2(net44),
    .B1(net28),
    .B2(net33),
    .X(_3178_));
 sky130_fd_sc_hd__nand3_1 _4070_ (.A(_3175_),
    .B(_3177_),
    .C(net195),
    .Y(_3179_));
 sky130_fd_sc_hd__a21o_1 _4071_ (.A1(_3177_),
    .A2(_3178_),
    .B1(_3175_),
    .X(_3180_));
 sky130_fd_sc_hd__a21o_1 _4072_ (.A1(_0270_),
    .A2(_1471_),
    .B1(_1460_),
    .X(_3181_));
 sky130_fd_sc_hd__and3_1 _4073_ (.A(_3179_),
    .B(_3180_),
    .C(_3181_),
    .X(_3182_));
 sky130_fd_sc_hd__a21oi_1 _4074_ (.A1(_3179_),
    .A2(_3180_),
    .B1(_3181_),
    .Y(_3183_));
 sky130_fd_sc_hd__nor2_1 _4075_ (.A(_3182_),
    .B(_3183_),
    .Y(_3184_));
 sky130_fd_sc_hd__xnor2_2 _4076_ (.A(_3174_),
    .B(_3184_),
    .Y(_3185_));
 sky130_fd_sc_hd__o21ai_2 _4077_ (.A1(_3168_),
    .A2(_1515_),
    .B1(_3185_),
    .Y(_3186_));
 sky130_fd_sc_hd__or3_1 _4078_ (.A(_3168_),
    .B(_1515_),
    .C(_3185_),
    .X(_3187_));
 sky130_fd_sc_hd__nand2_1 _4079_ (.A(_3186_),
    .B(_3187_),
    .Y(_3188_));
 sky130_fd_sc_hd__xnor2_2 _4080_ (.A(_1439_),
    .B(_3188_),
    .Y(_3189_));
 sky130_fd_sc_hd__xnor2_1 _4081_ (.A(_1548_),
    .B(_3189_),
    .Y(_3190_));
 sky130_fd_sc_hd__nor2_1 _4082_ (.A(_1657_),
    .B(_3189_),
    .Y(_3191_));
 sky130_fd_sc_hd__or4bb_4 _4083_ (.A(_0783_),
    .B(_1144_),
    .C_N(_1154_),
    .D_N(_1165_),
    .X(_3192_));
 sky130_fd_sc_hd__a211oi_1 _4084_ (.A1(_1657_),
    .A2(_3190_),
    .B1(_3191_),
    .C1(_3192_),
    .Y(_3193_));
 sky130_fd_sc_hd__a211o_2 _4085_ (.A1(_0652_),
    .A2(_2969_),
    .B1(_3167_),
    .C1(_3193_),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_4 _4086_ (.A(net123),
    .X(_3194_));
 sky130_fd_sc_hd__buf_4 _4087_ (.A(net61),
    .X(_3195_));
 sky130_fd_sc_hd__clkbuf_4 _4088_ (.A(_3195_),
    .X(_3196_));
 sky130_fd_sc_hd__buf_4 _4089_ (.A(_3196_),
    .X(_3197_));
 sky130_fd_sc_hd__buf_2 _4090_ (.A(_3197_),
    .X(_3198_));
 sky130_fd_sc_hd__and2_1 _4091_ (.A(_2412_),
    .B(_3198_),
    .X(_3199_));
 sky130_fd_sc_hd__o21a_2 _4092_ (.A1(_0980_),
    .A2(_0969_),
    .B1(_0870_),
    .X(_3200_));
 sky130_fd_sc_hd__and2_2 _4093_ (.A(_0063_),
    .B(_3161_),
    .X(_3201_));
 sky130_fd_sc_hd__or2_2 _4094_ (.A(_2401_),
    .B(_3198_),
    .X(_3202_));
 sky130_fd_sc_hd__o21ai_1 _4095_ (.A1(_1209_),
    .A2(_3199_),
    .B1(_3202_),
    .Y(_3203_));
 sky130_fd_sc_hd__buf_2 _4096_ (.A(_1220_),
    .X(_3204_));
 sky130_fd_sc_hd__o22a_1 _4097_ (.A1(_1187_),
    .A2(_3202_),
    .B1(_3203_),
    .B2(_3204_),
    .X(_3205_));
 sky130_fd_sc_hd__a221o_1 _4098_ (.A1(_3194_),
    .A2(_3199_),
    .B1(_3200_),
    .B2(_3201_),
    .C1(_3205_),
    .X(_3206_));
 sky130_fd_sc_hd__mux4_2 _4099_ (.A0(_2412_),
    .A1(_2346_),
    .A2(_1023_),
    .A3(_1034_),
    .S0(_0925_),
    .S1(_3131_),
    .X(_3207_));
 sky130_fd_sc_hd__mux2_1 _4100_ (.A0(_1045_),
    .A1(_1067_),
    .S(_0914_),
    .X(_3208_));
 sky130_fd_sc_hd__clkbuf_8 _4101_ (.A(_1384_),
    .X(_3209_));
 sky130_fd_sc_hd__or2b_2 _4102_ (.A(_0903_),
    .B_N(_3209_),
    .X(_3210_));
 sky130_fd_sc_hd__inv_2 _4103_ (.A(_3210_),
    .Y(_3211_));
 sky130_fd_sc_hd__mux2_1 _4104_ (.A0(_3208_),
    .A1(_3211_),
    .S(_3131_),
    .X(_3212_));
 sky130_fd_sc_hd__mux2_2 _4105_ (.A0(_3207_),
    .A1(_3212_),
    .S(_1100_),
    .X(_3213_));
 sky130_fd_sc_hd__nand2_1 _4106_ (.A(_2401_),
    .B(_3198_),
    .Y(_3214_));
 sky130_fd_sc_hd__nand2_2 _4107_ (.A(_3202_),
    .B(_3214_),
    .Y(_3215_));
 sky130_fd_sc_hd__a21oi_1 _4108_ (.A1(_3159_),
    .A2(_2991_),
    .B1(_2914_),
    .Y(_3216_));
 sky130_fd_sc_hd__xnor2_1 _4109_ (.A(_3215_),
    .B(_3216_),
    .Y(_3217_));
 sky130_fd_sc_hd__a32o_1 _4110_ (.A1(_0838_),
    .A2(_3126_),
    .A3(_3213_),
    .B1(_3217_),
    .B2(_2980_),
    .X(_3218_));
 sky130_fd_sc_hd__mux2_1 _4111_ (.A0(_2620_),
    .A1(_1920_),
    .S(_3131_),
    .X(_3219_));
 sky130_fd_sc_hd__mux2_1 _4112_ (.A0(_2795_),
    .A1(_2554_),
    .S(_3131_),
    .X(_3220_));
 sky130_fd_sc_hd__mux2_1 _4113_ (.A0(_2281_),
    .A1(_2729_),
    .S(_3131_),
    .X(_3221_));
 sky130_fd_sc_hd__mux2_1 _4114_ (.A0(_2467_),
    .A1(_2193_),
    .S(_3131_),
    .X(_3222_));
 sky130_fd_sc_hd__mux4_1 _4115_ (.A0(_3219_),
    .A1(_3220_),
    .A2(_3221_),
    .A3(_3222_),
    .S0(_1712_),
    .S1(_1723_),
    .X(_3223_));
 sky130_fd_sc_hd__mux2_1 _4116_ (.A0(_1832_),
    .A1(_2040_),
    .S(_0947_),
    .X(_3224_));
 sky130_fd_sc_hd__mux2_1 _4117_ (.A0(_1974_),
    .A1(_1788_),
    .S(_0947_),
    .X(_3225_));
 sky130_fd_sc_hd__mux2_1 _4118_ (.A0(_3224_),
    .A1(_3225_),
    .S(_1712_),
    .X(_3226_));
 sky130_fd_sc_hd__mux2_1 _4119_ (.A0(_2062_),
    .A1(_3226_),
    .S(_0587_),
    .X(_3227_));
 sky130_fd_sc_hd__or3b_2 _4120_ (.A(_3200_),
    .B(_3154_),
    .C_N(_3227_),
    .X(_3228_));
 sky130_fd_sc_hd__a2bb2o_1 _4121_ (.A1_N(_0063_),
    .A2_N(_3223_),
    .B1(_3228_),
    .B2(_3156_),
    .X(_3229_));
 sky130_fd_sc_hd__or2b_1 _4122_ (.A(_3218_),
    .B_N(_3229_),
    .X(_3230_));
 sky130_fd_sc_hd__nand3b_1 _4123_ (.A_N(_1439_),
    .B(_3186_),
    .C(_3187_),
    .Y(_3231_));
 sky130_fd_sc_hd__and3_1 _4124_ (.A(net1),
    .B(net60),
    .C(_3172_),
    .X(_3232_));
 sky130_fd_sc_hd__o211a_1 _4125_ (.A1(_3171_),
    .A2(_3232_),
    .B1(net1),
    .C1(_3197_),
    .X(_3233_));
 sky130_fd_sc_hd__a211oi_1 _4126_ (.A1(_0466_),
    .A2(_3197_),
    .B1(_3171_),
    .C1(_3232_),
    .Y(_3234_));
 sky130_fd_sc_hd__or2_1 _4127_ (.A(_3233_),
    .B(_3234_),
    .X(_3235_));
 sky130_fd_sc_hd__a22oi_2 _4128_ (.A1(_3169_),
    .A2(_1264_),
    .B1(_0314_),
    .B2(_0030_),
    .Y(_3236_));
 sky130_fd_sc_hd__and4_1 _4129_ (.A(net58),
    .B(net59),
    .C(_1264_),
    .D(_0314_),
    .X(_3237_));
 sky130_fd_sc_hd__nor2_1 _4130_ (.A(_3236_),
    .B(_3237_),
    .Y(_3238_));
 sky130_fd_sc_hd__nand2_1 _4131_ (.A(_0412_),
    .B(net60),
    .Y(_3239_));
 sky130_fd_sc_hd__xnor2_2 _4132_ (.A(_3238_),
    .B(_3239_),
    .Y(_3240_));
 sky130_fd_sc_hd__and2_1 _4133_ (.A(net55),
    .B(_0074_),
    .X(_3241_));
 sky130_fd_sc_hd__buf_6 _4134_ (.A(net33),
    .X(_3242_));
 sky130_fd_sc_hd__nand4_1 _4135_ (.A(_3242_),
    .B(net44),
    .C(net28),
    .D(net29),
    .Y(_3243_));
 sky130_fd_sc_hd__a22o_1 _4136_ (.A1(net44),
    .A2(net28),
    .B1(net29),
    .B2(net33),
    .X(_3244_));
 sky130_fd_sc_hd__nand3_1 _4137_ (.A(_3241_),
    .B(_3243_),
    .C(_3244_),
    .Y(_3245_));
 sky130_fd_sc_hd__a21o_1 _4138_ (.A1(_3243_),
    .A2(_3244_),
    .B1(_3241_),
    .X(_3246_));
 sky130_fd_sc_hd__a21bo_1 _4139_ (.A1(_3175_),
    .A2(_3178_),
    .B1_N(_3177_),
    .X(_3247_));
 sky130_fd_sc_hd__nand3_1 _4140_ (.A(_3245_),
    .B(_3246_),
    .C(_3247_),
    .Y(_3248_));
 sky130_fd_sc_hd__a21o_1 _4141_ (.A1(_3245_),
    .A2(_3246_),
    .B1(_3247_),
    .X(_3249_));
 sky130_fd_sc_hd__nand3_1 _4142_ (.A(_3240_),
    .B(_3248_),
    .C(_3249_),
    .Y(_3250_));
 sky130_fd_sc_hd__a21o_1 _4143_ (.A1(_3248_),
    .A2(_3249_),
    .B1(_3240_),
    .X(_3251_));
 sky130_fd_sc_hd__o21bai_1 _4144_ (.A1(_3174_),
    .A2(_3183_),
    .B1_N(_3182_),
    .Y(_3252_));
 sky130_fd_sc_hd__and3_1 _4145_ (.A(_3250_),
    .B(_3251_),
    .C(_3252_),
    .X(_3253_));
 sky130_fd_sc_hd__a21oi_1 _4146_ (.A1(_3250_),
    .A2(_3251_),
    .B1(_3252_),
    .Y(_3254_));
 sky130_fd_sc_hd__nor3_1 _4147_ (.A(_3235_),
    .B(_3253_),
    .C(_3254_),
    .Y(_3255_));
 sky130_fd_sc_hd__o21a_1 _4148_ (.A1(_3253_),
    .A2(_3254_),
    .B1(_3235_),
    .X(_3256_));
 sky130_fd_sc_hd__a211o_1 _4149_ (.A1(_3186_),
    .A2(_3231_),
    .B1(net159),
    .C1(_3256_),
    .X(_3257_));
 sky130_fd_sc_hd__o211ai_1 _4150_ (.A1(net160),
    .A2(_3256_),
    .B1(_3186_),
    .C1(_3231_),
    .Y(_3258_));
 sky130_fd_sc_hd__or4bb_2 _4151_ (.A(_1548_),
    .B(_3189_),
    .C_N(_3257_),
    .D_N(_3258_),
    .X(_3259_));
 sky130_fd_sc_hd__a2bb2o_1 _4152_ (.A1_N(_1548_),
    .A2_N(_3189_),
    .B1(_3257_),
    .B2(_3258_),
    .X(_3260_));
 sky130_fd_sc_hd__a21o_1 _4153_ (.A1(_3259_),
    .A2(_3260_),
    .B1(_3191_),
    .X(_3261_));
 sky130_fd_sc_hd__nand3_1 _4154_ (.A(_3191_),
    .B(net176),
    .C(_3260_),
    .Y(_3262_));
 sky130_fd_sc_hd__and2b_1 _4155_ (.A_N(_2903_),
    .B(_2335_),
    .X(_3263_));
 sky130_fd_sc_hd__a21o_1 _4156_ (.A1(_2936_),
    .A2(_2958_),
    .B1(_3263_),
    .X(_3264_));
 sky130_fd_sc_hd__or2_2 _4157_ (.A(_0630_),
    .B(_0641_),
    .X(_3265_));
 sky130_fd_sc_hd__a21oi_1 _4158_ (.A1(_3215_),
    .A2(_3264_),
    .B1(_3265_),
    .Y(_3266_));
 sky130_fd_sc_hd__o21a_1 _4159_ (.A1(_3215_),
    .A2(_3264_),
    .B1(_3266_),
    .X(_3267_));
 sky130_fd_sc_hd__a31o_1 _4160_ (.A1(_1668_),
    .A2(_3261_),
    .A3(_3262_),
    .B1(_3267_),
    .X(_3268_));
 sky130_fd_sc_hd__or3_1 _4161_ (.A(_3206_),
    .B(_3230_),
    .C(_3268_),
    .X(_3269_));
 sky130_fd_sc_hd__clkbuf_2 _4162_ (.A(_3269_),
    .X(net97));
 sky130_fd_sc_hd__buf_6 _4163_ (.A(net62),
    .X(_3270_));
 sky130_fd_sc_hd__clkbuf_4 _4164_ (.A(_3270_),
    .X(_3271_));
 sky130_fd_sc_hd__buf_4 _4165_ (.A(_3271_),
    .X(_3272_));
 sky130_fd_sc_hd__clkbuf_4 _4166_ (.A(_3272_),
    .X(_3273_));
 sky130_fd_sc_hd__and2_1 _4167_ (.A(_2456_),
    .B(_3273_),
    .X(_3274_));
 sky130_fd_sc_hd__nor2_1 _4168_ (.A(_2456_),
    .B(_3273_),
    .Y(_3275_));
 sky130_fd_sc_hd__or2_2 _4169_ (.A(_3274_),
    .B(_3275_),
    .X(_3276_));
 sky130_fd_sc_hd__and2b_1 _4170_ (.A_N(_3198_),
    .B(_2412_),
    .X(_3277_));
 sky130_fd_sc_hd__a21o_1 _4171_ (.A1(_3215_),
    .A2(_3264_),
    .B1(_3277_),
    .X(_3278_));
 sky130_fd_sc_hd__nand2_1 _4172_ (.A(_3276_),
    .B(_3278_),
    .Y(_3279_));
 sky130_fd_sc_hd__o21a_1 _4173_ (.A1(_3276_),
    .A2(_3278_),
    .B1(_0652_),
    .X(_3280_));
 sky130_fd_sc_hd__a21o_1 _4174_ (.A1(_3202_),
    .A2(_3216_),
    .B1(_3199_),
    .X(_3281_));
 sky130_fd_sc_hd__xnor2_1 _4175_ (.A(_3276_),
    .B(_3281_),
    .Y(_3282_));
 sky130_fd_sc_hd__mux4_2 _4176_ (.A0(_3139_),
    .A1(_2412_),
    .A2(_2346_),
    .A3(_1023_),
    .S0(_0925_),
    .S1(_0969_),
    .X(_3283_));
 sky130_fd_sc_hd__mux4_2 _4177_ (.A0(_1034_),
    .A1(_1045_),
    .A2(_1067_),
    .A3(_3209_),
    .S0(_0914_),
    .S1(_0958_),
    .X(_3284_));
 sky130_fd_sc_hd__mux2_2 _4178_ (.A0(_3283_),
    .A1(_3284_),
    .S(_1100_),
    .X(_3285_));
 sky130_fd_sc_hd__o21ba_1 _4179_ (.A1(_1209_),
    .A2(_3274_),
    .B1_N(_3204_),
    .X(_3286_));
 sky130_fd_sc_hd__nor2_1 _4180_ (.A(_3275_),
    .B(_3286_),
    .Y(_3287_));
 sky130_fd_sc_hd__a221o_1 _4181_ (.A1(net123),
    .A2(_3274_),
    .B1(_3275_),
    .B2(_1187_),
    .C1(_3162_),
    .X(_3288_));
 sky130_fd_sc_hd__a311o_1 _4182_ (.A1(_0838_),
    .A2(_3126_),
    .A3(_3285_),
    .B1(_3287_),
    .C1(_3288_),
    .X(_3289_));
 sky130_fd_sc_hd__nor2_1 _4183_ (.A(_0947_),
    .B(_3147_),
    .Y(_3290_));
 sky130_fd_sc_hd__a21oi_1 _4184_ (.A1(_0947_),
    .A2(_3143_),
    .B1(_3290_),
    .Y(_3291_));
 sky130_fd_sc_hd__mux2_1 _4185_ (.A0(_3150_),
    .A1(_3146_),
    .S(_0521_),
    .X(_3292_));
 sky130_fd_sc_hd__mux2_1 _4186_ (.A0(_3291_),
    .A1(_3292_),
    .S(_1712_),
    .X(_3293_));
 sky130_fd_sc_hd__nor2_1 _4187_ (.A(_3108_),
    .B(_3293_),
    .Y(_3294_));
 sky130_fd_sc_hd__a2111o_1 _4188_ (.A1(_3108_),
    .A2(_3144_),
    .B1(_3200_),
    .C1(_3294_),
    .D1(_3154_),
    .X(_3295_));
 sky130_fd_sc_hd__mux2_1 _4189_ (.A0(_3130_),
    .A1(_3149_),
    .S(_0936_),
    .X(_3296_));
 sky130_fd_sc_hd__mux2_1 _4190_ (.A0(_3135_),
    .A1(_2510_),
    .S(_0903_),
    .X(_3297_));
 sky130_fd_sc_hd__mux2_1 _4191_ (.A0(_3297_),
    .A1(_3129_),
    .S(_0958_),
    .X(_3298_));
 sky130_fd_sc_hd__mux4_1 _4192_ (.A0(_3137_),
    .A1(_2675_),
    .A2(_3133_),
    .A3(_2762_),
    .S0(_0903_),
    .S1(_0958_),
    .X(_3299_));
 sky130_fd_sc_hd__mux4_1 _4193_ (.A0(_3139_),
    .A1(_2138_),
    .A2(_2182_),
    .A3(_2237_),
    .S0(_0903_),
    .S1(_0958_),
    .X(_3300_));
 sky130_fd_sc_hd__clkbuf_4 _4194_ (.A(_1723_),
    .X(_3301_));
 sky130_fd_sc_hd__mux4_1 _4195_ (.A0(_3296_),
    .A1(_3298_),
    .A2(_3299_),
    .A3(_3300_),
    .S0(_3077_),
    .S1(_3301_),
    .X(_3302_));
 sky130_fd_sc_hd__o2bb2a_1 _4196_ (.A1_N(_3156_),
    .A2_N(_3295_),
    .B1(_3302_),
    .B2(_3127_),
    .X(_3303_));
 sky130_fd_sc_hd__a211o_1 _4197_ (.A1(_2980_),
    .A2(_3282_),
    .B1(_3289_),
    .C1(_3303_),
    .X(_3304_));
 sky130_fd_sc_hd__buf_4 _4198_ (.A(_1668_),
    .X(_3305_));
 sky130_fd_sc_hd__o21ba_1 _4199_ (.A1(_3236_),
    .A2(_3239_),
    .B1_N(_3237_),
    .X(_3306_));
 sky130_fd_sc_hd__a22oi_2 _4200_ (.A1(_0434_),
    .A2(_3196_),
    .B1(_3272_),
    .B2(net1),
    .Y(_3307_));
 sky130_fd_sc_hd__and4_1 _4201_ (.A(net163),
    .B(net1),
    .C(_3196_),
    .D(_3271_),
    .X(_3308_));
 sky130_fd_sc_hd__nor2_1 _4202_ (.A(_3307_),
    .B(_3308_),
    .Y(_3309_));
 sky130_fd_sc_hd__xnor2_2 _4203_ (.A(_3306_),
    .B(_3309_),
    .Y(_3310_));
 sky130_fd_sc_hd__nand2_1 _4204_ (.A(_0324_),
    .B(net60),
    .Y(_3311_));
 sky130_fd_sc_hd__and4_1 _4205_ (.A(net58),
    .B(net59),
    .C(net27),
    .D(net26),
    .X(_3312_));
 sky130_fd_sc_hd__a22o_1 _4206_ (.A1(net58),
    .A2(_0074_),
    .B1(net26),
    .B2(net59),
    .X(_3313_));
 sky130_fd_sc_hd__and2b_1 _4207_ (.A_N(_3312_),
    .B(_3313_),
    .X(_3314_));
 sky130_fd_sc_hd__xnor2_2 _4208_ (.A(_3311_),
    .B(_3314_),
    .Y(_3315_));
 sky130_fd_sc_hd__and2_1 _4209_ (.A(net55),
    .B(net28),
    .X(_3316_));
 sky130_fd_sc_hd__nand4_2 _4210_ (.A(_3242_),
    .B(_3176_),
    .C(net29),
    .D(net30),
    .Y(_3317_));
 sky130_fd_sc_hd__a22o_1 _4211_ (.A1(net44),
    .A2(net29),
    .B1(net30),
    .B2(net33),
    .X(_3318_));
 sky130_fd_sc_hd__nand3_1 _4212_ (.A(_3316_),
    .B(_3317_),
    .C(_3318_),
    .Y(_3319_));
 sky130_fd_sc_hd__a21o_1 _4213_ (.A1(_3317_),
    .A2(_3318_),
    .B1(_3316_),
    .X(_3320_));
 sky130_fd_sc_hd__a21bo_1 _4214_ (.A1(_3241_),
    .A2(_3244_),
    .B1_N(_3243_),
    .X(_3321_));
 sky130_fd_sc_hd__nand3_1 _4215_ (.A(_3319_),
    .B(_3320_),
    .C(_3321_),
    .Y(_3322_));
 sky130_fd_sc_hd__a21o_1 _4216_ (.A1(_3319_),
    .A2(_3320_),
    .B1(_3321_),
    .X(_3323_));
 sky130_fd_sc_hd__nand3_1 _4217_ (.A(_3315_),
    .B(_3322_),
    .C(_3323_),
    .Y(_3324_));
 sky130_fd_sc_hd__a21o_1 _4218_ (.A1(_3322_),
    .A2(_3323_),
    .B1(_3315_),
    .X(_3325_));
 sky130_fd_sc_hd__a21bo_1 _4219_ (.A1(_3240_),
    .A2(_3249_),
    .B1_N(_3248_),
    .X(_3326_));
 sky130_fd_sc_hd__nand3_2 _4220_ (.A(_3324_),
    .B(_3325_),
    .C(_3326_),
    .Y(_3327_));
 sky130_fd_sc_hd__a21o_1 _4221_ (.A1(_3324_),
    .A2(_3325_),
    .B1(_3326_),
    .X(_3328_));
 sky130_fd_sc_hd__nand3_2 _4222_ (.A(_3310_),
    .B(_3327_),
    .C(_3328_),
    .Y(_3329_));
 sky130_fd_sc_hd__a21o_1 _4223_ (.A1(_3327_),
    .A2(_3328_),
    .B1(_3310_),
    .X(_3330_));
 sky130_fd_sc_hd__o211a_1 _4224_ (.A1(_3253_),
    .A2(_3255_),
    .B1(_3329_),
    .C1(_3330_),
    .X(_3331_));
 sky130_fd_sc_hd__a211o_1 _4225_ (.A1(_3329_),
    .A2(_3330_),
    .B1(_3253_),
    .C1(_3255_),
    .X(_3332_));
 sky130_fd_sc_hd__and2b_1 _4226_ (.A_N(_3331_),
    .B(_3332_),
    .X(_3333_));
 sky130_fd_sc_hd__xnor2_2 _4227_ (.A(net193),
    .B(_3333_),
    .Y(_3334_));
 sky130_fd_sc_hd__nand2_1 _4228_ (.A(net145),
    .B(_3259_),
    .Y(_3335_));
 sky130_fd_sc_hd__xor2_1 _4229_ (.A(net192),
    .B(_3335_),
    .X(_3336_));
 sky130_fd_sc_hd__nand2_1 _4230_ (.A(_3262_),
    .B(_3336_),
    .Y(_3337_));
 sky130_fd_sc_hd__or2_1 _4231_ (.A(_3262_),
    .B(_3336_),
    .X(_3338_));
 sky130_fd_sc_hd__and3_1 _4232_ (.A(_3305_),
    .B(_3337_),
    .C(_3338_),
    .X(_3339_));
 sky130_fd_sc_hd__a211o_4 _4233_ (.A1(_3279_),
    .A2(_3280_),
    .B1(_3304_),
    .C1(_3339_),
    .X(net98));
 sky130_fd_sc_hd__or3_2 _4234_ (.A(_3306_),
    .B(_3307_),
    .C(_3308_),
    .X(_3340_));
 sky130_fd_sc_hd__inv_2 _4235_ (.A(_3308_),
    .Y(_3341_));
 sky130_fd_sc_hd__a31o_1 _4236_ (.A1(_0324_),
    .A2(net60),
    .A3(_3313_),
    .B1(_3312_),
    .X(_3342_));
 sky130_fd_sc_hd__buf_2 _4237_ (.A(net63),
    .X(_3343_));
 sky130_fd_sc_hd__a22oi_1 _4238_ (.A1(net23),
    .A2(net61),
    .B1(_3270_),
    .B2(_0412_),
    .Y(_3344_));
 sky130_fd_sc_hd__and4_1 _4239_ (.A(net23),
    .B(net12),
    .C(net61),
    .D(net62),
    .X(_3345_));
 sky130_fd_sc_hd__o2bb2a_1 _4240_ (.A1_N(net1),
    .A2_N(_3343_),
    .B1(_3344_),
    .B2(_3345_),
    .X(_3346_));
 sky130_fd_sc_hd__and4bb_1 _4241_ (.A_N(_3344_),
    .B_N(_3345_),
    .C(net1),
    .D(net63),
    .X(_3347_));
 sky130_fd_sc_hd__or2_2 _4242_ (.A(_3346_),
    .B(_3347_),
    .X(_3348_));
 sky130_fd_sc_hd__xor2_2 _4243_ (.A(_3342_),
    .B(_3348_),
    .X(_3349_));
 sky130_fd_sc_hd__xnor2_1 _4244_ (.A(_3341_),
    .B(_3349_),
    .Y(_3350_));
 sky130_fd_sc_hd__nand2_1 _4245_ (.A(_0194_),
    .B(net60),
    .Y(_3351_));
 sky130_fd_sc_hd__clkbuf_4 _4246_ (.A(net58),
    .X(_3352_));
 sky130_fd_sc_hd__and3_1 _4247_ (.A(net59),
    .B(_0074_),
    .C(net28),
    .X(_3353_));
 sky130_fd_sc_hd__a22o_1 _4248_ (.A1(net59),
    .A2(_0074_),
    .B1(net28),
    .B2(net58),
    .X(_3354_));
 sky130_fd_sc_hd__a21bo_1 _4249_ (.A1(_3352_),
    .A2(_3353_),
    .B1_N(_3354_),
    .X(_3355_));
 sky130_fd_sc_hd__xor2_2 _4250_ (.A(_3351_),
    .B(_3355_),
    .X(_3356_));
 sky130_fd_sc_hd__and2_1 _4251_ (.A(net55),
    .B(net29),
    .X(_3357_));
 sky130_fd_sc_hd__nand4_2 _4252_ (.A(_3242_),
    .B(_3176_),
    .C(net30),
    .D(net31),
    .Y(_3358_));
 sky130_fd_sc_hd__a22o_1 _4253_ (.A1(net44),
    .A2(net30),
    .B1(net31),
    .B2(net33),
    .X(_3359_));
 sky130_fd_sc_hd__nand3_1 _4254_ (.A(_3357_),
    .B(_3358_),
    .C(_3359_),
    .Y(_3360_));
 sky130_fd_sc_hd__a21o_1 _4255_ (.A1(_3358_),
    .A2(_3359_),
    .B1(_3357_),
    .X(_3361_));
 sky130_fd_sc_hd__a21bo_1 _4256_ (.A1(_3316_),
    .A2(_3318_),
    .B1_N(_3317_),
    .X(_3362_));
 sky130_fd_sc_hd__nand3_1 _4257_ (.A(_3360_),
    .B(_3361_),
    .C(_3362_),
    .Y(_3363_));
 sky130_fd_sc_hd__a21o_1 _4258_ (.A1(_3360_),
    .A2(_3361_),
    .B1(_3362_),
    .X(_3364_));
 sky130_fd_sc_hd__nand3_1 _4259_ (.A(_3356_),
    .B(_3363_),
    .C(_3364_),
    .Y(_3365_));
 sky130_fd_sc_hd__a21o_1 _4260_ (.A1(_3363_),
    .A2(_3364_),
    .B1(_3356_),
    .X(_3366_));
 sky130_fd_sc_hd__a21bo_1 _4261_ (.A1(_3315_),
    .A2(_3323_),
    .B1_N(_3322_),
    .X(_3367_));
 sky130_fd_sc_hd__and3_2 _4262_ (.A(_3365_),
    .B(_3366_),
    .C(_3367_),
    .X(_3368_));
 sky130_fd_sc_hd__a21oi_1 _4263_ (.A1(_3365_),
    .A2(_3366_),
    .B1(_3367_),
    .Y(_3369_));
 sky130_fd_sc_hd__nor3_1 _4264_ (.A(_3350_),
    .B(_3368_),
    .C(_3369_),
    .Y(_3370_));
 sky130_fd_sc_hd__o21a_1 _4265_ (.A1(_3368_),
    .A2(_3369_),
    .B1(_3350_),
    .X(_3371_));
 sky130_fd_sc_hd__a211oi_2 _4266_ (.A1(_3327_),
    .A2(_3329_),
    .B1(_3370_),
    .C1(net184),
    .Y(_3372_));
 sky130_fd_sc_hd__o211a_1 _4267_ (.A1(_3370_),
    .A2(_3371_),
    .B1(_3327_),
    .C1(_3329_),
    .X(_3373_));
 sky130_fd_sc_hd__or3_1 _4268_ (.A(_3340_),
    .B(_3372_),
    .C(_3373_),
    .X(_3374_));
 sky130_fd_sc_hd__o21ai_2 _4269_ (.A1(_3372_),
    .A2(_3373_),
    .B1(_3340_),
    .Y(_3375_));
 sky130_fd_sc_hd__a21o_1 _4270_ (.A1(net193),
    .A2(_3332_),
    .B1(_3331_),
    .X(_3376_));
 sky130_fd_sc_hd__and3_1 _4271_ (.A(_3374_),
    .B(_3375_),
    .C(_3376_),
    .X(_3377_));
 sky130_fd_sc_hd__a21oi_2 _4272_ (.A1(net186),
    .A2(_3375_),
    .B1(net196),
    .Y(_3378_));
 sky130_fd_sc_hd__or4_1 _4273_ (.A(_3257_),
    .B(_3334_),
    .C(_3377_),
    .D(_3378_),
    .X(_3379_));
 sky130_fd_sc_hd__o22ai_1 _4274_ (.A1(net147),
    .A2(_3334_),
    .B1(_3377_),
    .B2(_3378_),
    .Y(_3380_));
 sky130_fd_sc_hd__or4bb_2 _4275_ (.A(_3259_),
    .B(net192),
    .C_N(_3379_),
    .D_N(_3380_),
    .X(_3381_));
 sky130_fd_sc_hd__a2bb2o_1 _4276_ (.A1_N(_3259_),
    .A2_N(net192),
    .B1(net188),
    .B2(_3380_),
    .X(_3382_));
 sky130_fd_sc_hd__a21bo_1 _4277_ (.A1(_3381_),
    .A2(_3382_),
    .B1_N(_3338_),
    .X(_3383_));
 sky130_fd_sc_hd__or4bb_1 _4278_ (.A(_3262_),
    .B(_3336_),
    .C_N(_3381_),
    .D_N(_3382_),
    .X(_3384_));
 sky130_fd_sc_hd__clkbuf_4 _4279_ (.A(_3343_),
    .X(_3385_));
 sky130_fd_sc_hd__clkbuf_4 _4280_ (.A(_3385_),
    .X(_3386_));
 sky130_fd_sc_hd__nor2_1 _4281_ (.A(_2127_),
    .B(_3386_),
    .Y(_3387_));
 sky130_fd_sc_hd__and2_4 _4282_ (.A(net31),
    .B(net63),
    .X(_3388_));
 sky130_fd_sc_hd__or2_2 _4283_ (.A(_3387_),
    .B(_3388_),
    .X(_3389_));
 sky130_fd_sc_hd__and2b_1 _4284_ (.A_N(_3273_),
    .B(_3139_),
    .X(_3390_));
 sky130_fd_sc_hd__a21o_1 _4285_ (.A1(_3276_),
    .A2(_3278_),
    .B1(_3390_),
    .X(_3391_));
 sky130_fd_sc_hd__or2_1 _4286_ (.A(_3389_),
    .B(_3391_),
    .X(_3392_));
 sky130_fd_sc_hd__nand2_1 _4287_ (.A(_3389_),
    .B(_3391_),
    .Y(_3393_));
 sky130_fd_sc_hd__o211a_1 _4288_ (.A1(_2456_),
    .A2(_3273_),
    .B1(_2401_),
    .C1(_3198_),
    .X(_3394_));
 sky130_fd_sc_hd__nor2_1 _4289_ (.A(_3274_),
    .B(_3394_),
    .Y(_3395_));
 sky130_fd_sc_hd__a2111o_1 _4290_ (.A1(_3159_),
    .A2(_2991_),
    .B1(_3215_),
    .C1(_3276_),
    .D1(_2914_),
    .X(_3396_));
 sky130_fd_sc_hd__and2_1 _4291_ (.A(_3395_),
    .B(_3396_),
    .X(_3397_));
 sky130_fd_sc_hd__nand2_1 _4292_ (.A(_3389_),
    .B(_3397_),
    .Y(_3398_));
 sky130_fd_sc_hd__o21a_1 _4293_ (.A1(_3389_),
    .A2(_3397_),
    .B1(_2980_),
    .X(_3399_));
 sky130_fd_sc_hd__mux2_1 _4294_ (.A0(_2292_),
    .A1(_2806_),
    .S(_1100_),
    .X(_3400_));
 sky130_fd_sc_hd__mux2_1 _4295_ (.A0(_1985_),
    .A1(_2631_),
    .S(_1712_),
    .X(_3401_));
 sky130_fd_sc_hd__mux2_1 _4296_ (.A0(_3400_),
    .A1(_3401_),
    .S(_0870_),
    .X(_3402_));
 sky130_fd_sc_hd__mux2_1 _4297_ (.A0(_2073_),
    .A1(_1843_),
    .S(_1712_),
    .X(_3403_));
 sky130_fd_sc_hd__nand2_1 _4298_ (.A(_1723_),
    .B(_3403_),
    .Y(_3404_));
 sky130_fd_sc_hd__nand2_1 _4299_ (.A(_3127_),
    .B(_3404_),
    .Y(_3405_));
 sky130_fd_sc_hd__o211a_1 _4300_ (.A1(_3127_),
    .A2(_3402_),
    .B1(_3405_),
    .C1(_1701_),
    .X(_3406_));
 sky130_fd_sc_hd__mux4_2 _4301_ (.A0(_2138_),
    .A1(_3139_),
    .A2(_2412_),
    .A3(_2346_),
    .S0(_0914_),
    .S1(_3131_),
    .X(_3407_));
 sky130_fd_sc_hd__nand2_1 _4302_ (.A(_3077_),
    .B(_3407_),
    .Y(_3408_));
 sky130_fd_sc_hd__o211a_1 _4303_ (.A1(_3077_),
    .A2(_1089_),
    .B1(_3408_),
    .C1(_1723_),
    .X(_3409_));
 sky130_fd_sc_hd__a211o_1 _4304_ (.A1(_3108_),
    .A2(_3210_),
    .B1(_3409_),
    .C1(_3200_),
    .X(_3410_));
 sky130_fd_sc_hd__nor2_1 _4305_ (.A(_0860_),
    .B(_3410_),
    .Y(_3411_));
 sky130_fd_sc_hd__o21ba_1 _4306_ (.A1(_1209_),
    .A2(_3388_),
    .B1_N(_3204_),
    .X(_3412_));
 sky130_fd_sc_hd__nor2_1 _4307_ (.A(_3387_),
    .B(_3412_),
    .Y(_3413_));
 sky130_fd_sc_hd__clkbuf_4 _4308_ (.A(_1187_),
    .X(_3414_));
 sky130_fd_sc_hd__a221o_1 _4309_ (.A1(_3414_),
    .A2(_3387_),
    .B1(_3388_),
    .B2(net123),
    .C1(_3162_),
    .X(_3415_));
 sky130_fd_sc_hd__or4_1 _4310_ (.A(_3406_),
    .B(_3411_),
    .C(_3413_),
    .D(_3415_),
    .X(_3416_));
 sky130_fd_sc_hd__a21o_1 _4311_ (.A1(_3398_),
    .A2(_3399_),
    .B1(_3416_),
    .X(_3417_));
 sky130_fd_sc_hd__a31o_1 _4312_ (.A1(_0652_),
    .A2(_3392_),
    .A3(_3393_),
    .B1(_3417_),
    .X(_3418_));
 sky130_fd_sc_hd__a31o_2 _4313_ (.A1(_3305_),
    .A2(_3383_),
    .A3(_3384_),
    .B1(_3418_),
    .X(net99));
 sky130_fd_sc_hd__nor3_1 _4314_ (.A(_3340_),
    .B(_3372_),
    .C(_3373_),
    .Y(_3419_));
 sky130_fd_sc_hd__or2b_1 _4315_ (.A(_3348_),
    .B_N(_3342_),
    .X(_3420_));
 sky130_fd_sc_hd__o21ai_2 _4316_ (.A1(_3341_),
    .A2(_3349_),
    .B1(_3420_),
    .Y(_3421_));
 sky130_fd_sc_hd__clkbuf_4 _4317_ (.A(net64),
    .X(_3422_));
 sky130_fd_sc_hd__clkbuf_4 _4318_ (.A(_3422_),
    .X(_3423_));
 sky130_fd_sc_hd__clkbuf_4 _4319_ (.A(_3423_),
    .X(_3424_));
 sky130_fd_sc_hd__clkbuf_4 _4320_ (.A(_3424_),
    .X(_3425_));
 sky130_fd_sc_hd__nand2_1 _4321_ (.A(_1002_),
    .B(_3425_),
    .Y(_3426_));
 sky130_fd_sc_hd__xnor2_2 _4322_ (.A(_3421_),
    .B(_3426_),
    .Y(_3427_));
 sky130_fd_sc_hd__or2_2 _4323_ (.A(_3345_),
    .B(_3347_),
    .X(_3428_));
 sky130_fd_sc_hd__a32o_1 _4324_ (.A1(_0205_),
    .A2(_2892_),
    .A3(_3354_),
    .B1(_3353_),
    .B2(_0172_),
    .X(_3429_));
 sky130_fd_sc_hd__clkbuf_4 _4325_ (.A(_3343_),
    .X(_3430_));
 sky130_fd_sc_hd__buf_4 _4326_ (.A(_3270_),
    .X(_3431_));
 sky130_fd_sc_hd__a22o_1 _4327_ (.A1(_1264_),
    .A2(net61),
    .B1(_3431_),
    .B2(_0314_),
    .X(_3432_));
 sky130_fd_sc_hd__clkbuf_4 _4328_ (.A(net61),
    .X(_3433_));
 sky130_fd_sc_hd__nand4_1 _4329_ (.A(_0194_),
    .B(_0314_),
    .C(_3433_),
    .D(_3431_),
    .Y(_3434_));
 sky130_fd_sc_hd__a22oi_1 _4330_ (.A1(_0423_),
    .A2(_3430_),
    .B1(_3432_),
    .B2(_3434_),
    .Y(_3435_));
 sky130_fd_sc_hd__and4_1 _4331_ (.A(net163),
    .B(_3343_),
    .C(_3432_),
    .D(_3434_),
    .X(_3436_));
 sky130_fd_sc_hd__or2_1 _4332_ (.A(_3435_),
    .B(_3436_),
    .X(_3437_));
 sky130_fd_sc_hd__xnor2_1 _4333_ (.A(_3429_),
    .B(_3437_),
    .Y(_3438_));
 sky130_fd_sc_hd__xor2_2 _4334_ (.A(_3428_),
    .B(_3438_),
    .X(_3439_));
 sky130_fd_sc_hd__clkbuf_4 _4335_ (.A(net194),
    .X(_3440_));
 sky130_fd_sc_hd__nand2_1 _4336_ (.A(_3440_),
    .B(_2881_),
    .Y(_3441_));
 sky130_fd_sc_hd__buf_4 _4337_ (.A(net29),
    .X(_3442_));
 sky130_fd_sc_hd__and3_1 _4338_ (.A(_3169_),
    .B(net191),
    .C(_2302_),
    .X(_3443_));
 sky130_fd_sc_hd__a22o_1 _4339_ (.A1(_0030_),
    .A2(_2302_),
    .B1(_2368_),
    .B2(_3169_),
    .X(_3444_));
 sky130_fd_sc_hd__a21bo_1 _4340_ (.A1(_3442_),
    .A2(_3443_),
    .B1_N(_3444_),
    .X(_3445_));
 sky130_fd_sc_hd__xor2_2 _4341_ (.A(_3441_),
    .B(_3445_),
    .X(_3446_));
 sky130_fd_sc_hd__and2_1 _4342_ (.A(_0292_),
    .B(_2423_),
    .X(_3447_));
 sky130_fd_sc_hd__buf_6 _4343_ (.A(_3176_),
    .X(_3448_));
 sky130_fd_sc_hd__buf_4 _4344_ (.A(_3242_),
    .X(_3449_));
 sky130_fd_sc_hd__a22o_1 _4345_ (.A1(_3448_),
    .A2(net31),
    .B1(net32),
    .B2(_3449_),
    .X(_3450_));
 sky130_fd_sc_hd__buf_4 _4346_ (.A(_3242_),
    .X(_3451_));
 sky130_fd_sc_hd__buf_4 _4347_ (.A(_3176_),
    .X(_3452_));
 sky130_fd_sc_hd__nand4_2 _4348_ (.A(_3451_),
    .B(_3452_),
    .C(_2106_),
    .D(_2149_),
    .Y(_3453_));
 sky130_fd_sc_hd__nand3_1 _4349_ (.A(_3447_),
    .B(_3450_),
    .C(_3453_),
    .Y(_3454_));
 sky130_fd_sc_hd__a21o_1 _4350_ (.A1(_3450_),
    .A2(_3453_),
    .B1(_3447_),
    .X(_3455_));
 sky130_fd_sc_hd__a21bo_1 _4351_ (.A1(_3357_),
    .A2(_3359_),
    .B1_N(_3358_),
    .X(_3456_));
 sky130_fd_sc_hd__nand3_1 _4352_ (.A(_3454_),
    .B(_3455_),
    .C(_3456_),
    .Y(_3457_));
 sky130_fd_sc_hd__a21o_1 _4353_ (.A1(_3454_),
    .A2(_3455_),
    .B1(_3456_),
    .X(_3458_));
 sky130_fd_sc_hd__nand3_2 _4354_ (.A(_3446_),
    .B(_3457_),
    .C(_3458_),
    .Y(_3459_));
 sky130_fd_sc_hd__a21o_1 _4355_ (.A1(_3457_),
    .A2(_3458_),
    .B1(_3446_),
    .X(_3460_));
 sky130_fd_sc_hd__a21bo_1 _4356_ (.A1(_3356_),
    .A2(_3364_),
    .B1_N(_3363_),
    .X(_3461_));
 sky130_fd_sc_hd__nand3_4 _4357_ (.A(_3459_),
    .B(_3460_),
    .C(_3461_),
    .Y(_3462_));
 sky130_fd_sc_hd__a21o_1 _4358_ (.A1(_3459_),
    .A2(_3460_),
    .B1(_3461_),
    .X(_3463_));
 sky130_fd_sc_hd__nand3_4 _4359_ (.A(_3439_),
    .B(_3462_),
    .C(_3463_),
    .Y(_3464_));
 sky130_fd_sc_hd__a21o_1 _4360_ (.A1(_3462_),
    .A2(_3463_),
    .B1(_3439_),
    .X(_3465_));
 sky130_fd_sc_hd__o211ai_4 _4361_ (.A1(_3368_),
    .A2(net122),
    .B1(_3464_),
    .C1(_3465_),
    .Y(_3466_));
 sky130_fd_sc_hd__a211o_1 _4362_ (.A1(_3464_),
    .A2(_3465_),
    .B1(_3368_),
    .C1(net122),
    .X(_3467_));
 sky130_fd_sc_hd__nand3_2 _4363_ (.A(_3427_),
    .B(_3466_),
    .C(_3467_),
    .Y(_3468_));
 sky130_fd_sc_hd__a21o_1 _4364_ (.A1(_3466_),
    .A2(_3467_),
    .B1(_3427_),
    .X(_3469_));
 sky130_fd_sc_hd__o211a_1 _4365_ (.A1(net183),
    .A2(_3419_),
    .B1(_3468_),
    .C1(_3469_),
    .X(_3470_));
 sky130_fd_sc_hd__a211o_1 _4366_ (.A1(_3468_),
    .A2(_3469_),
    .B1(net183),
    .C1(_3419_),
    .X(_3471_));
 sky130_fd_sc_hd__or2b_1 _4367_ (.A(_3470_),
    .B_N(_3471_),
    .X(_3472_));
 sky130_fd_sc_hd__nand3_1 _4368_ (.A(_3374_),
    .B(_3375_),
    .C(_3376_),
    .Y(_3473_));
 sky130_fd_sc_hd__o31ai_1 _4369_ (.A1(net146),
    .A2(_3334_),
    .A3(_3378_),
    .B1(_3473_),
    .Y(_3474_));
 sky130_fd_sc_hd__xor2_1 _4370_ (.A(_3472_),
    .B(_3474_),
    .X(_3475_));
 sky130_fd_sc_hd__nor2_1 _4371_ (.A(_3381_),
    .B(_3475_),
    .Y(_3476_));
 sky130_fd_sc_hd__and2_1 _4372_ (.A(_3381_),
    .B(_3475_),
    .X(_3477_));
 sky130_fd_sc_hd__o21ai_1 _4373_ (.A1(_3476_),
    .A2(_3477_),
    .B1(_3384_),
    .Y(_3478_));
 sky130_fd_sc_hd__or2_1 _4374_ (.A(_3384_),
    .B(_3475_),
    .X(_3479_));
 sky130_fd_sc_hd__and2_1 _4375_ (.A(_2171_),
    .B(_3425_),
    .X(_3480_));
 sky130_fd_sc_hd__nor2_1 _4376_ (.A(_2171_),
    .B(_3425_),
    .Y(_3481_));
 sky130_fd_sc_hd__or2_2 _4377_ (.A(_3480_),
    .B(_3481_),
    .X(_3482_));
 sky130_fd_sc_hd__o21ba_1 _4378_ (.A1(_3387_),
    .A2(_3397_),
    .B1_N(_3388_),
    .X(_3483_));
 sky130_fd_sc_hd__or2_1 _4379_ (.A(_3482_),
    .B(_3483_),
    .X(_3484_));
 sky130_fd_sc_hd__nand2_1 _4380_ (.A(_3482_),
    .B(_3483_),
    .Y(_3485_));
 sky130_fd_sc_hd__clkbuf_4 _4381_ (.A(_3108_),
    .X(_3486_));
 sky130_fd_sc_hd__and3_1 _4382_ (.A(_1100_),
    .B(_0925_),
    .C(_0969_),
    .X(_3487_));
 sky130_fd_sc_hd__o21a_1 _4383_ (.A1(_3486_),
    .A2(_3487_),
    .B1(_3201_),
    .X(_3488_));
 sky130_fd_sc_hd__a221o_1 _4384_ (.A1(_3194_),
    .A2(_3480_),
    .B1(_3481_),
    .B2(_3414_),
    .C1(_3488_),
    .X(_3489_));
 sky130_fd_sc_hd__clkbuf_4 _4385_ (.A(_1100_),
    .X(_3490_));
 sky130_fd_sc_hd__mux4_1 _4386_ (.A0(_3132_),
    .A1(_3138_),
    .A2(_3151_),
    .A3(_3136_),
    .S0(_1723_),
    .S1(_3490_),
    .X(_3491_));
 sky130_fd_sc_hd__nor2_1 _4387_ (.A(_0980_),
    .B(_3148_),
    .Y(_3492_));
 sky130_fd_sc_hd__a211o_1 _4388_ (.A1(_3490_),
    .A2(_3145_),
    .B1(_3492_),
    .C1(_3108_),
    .X(_3493_));
 sky130_fd_sc_hd__nand2_1 _4389_ (.A(_3127_),
    .B(_3493_),
    .Y(_3494_));
 sky130_fd_sc_hd__o211a_1 _4390_ (.A1(_3127_),
    .A2(_3491_),
    .B1(_3494_),
    .C1(_1701_),
    .X(_3495_));
 sky130_fd_sc_hd__and2b_1 _4391_ (.A_N(_3386_),
    .B(_2138_),
    .X(_3496_));
 sky130_fd_sc_hd__a21o_1 _4392_ (.A1(_3389_),
    .A2(_3391_),
    .B1(_3496_),
    .X(_3497_));
 sky130_fd_sc_hd__a21oi_1 _4393_ (.A1(_3482_),
    .A2(_3497_),
    .B1(_3265_),
    .Y(_3498_));
 sky130_fd_sc_hd__o21a_1 _4394_ (.A1(_3482_),
    .A2(_3497_),
    .B1(_3498_),
    .X(_3499_));
 sky130_fd_sc_hd__mux4_2 _4395_ (.A0(_2182_),
    .A1(_2138_),
    .A2(_3139_),
    .A3(_2412_),
    .S0(_0914_),
    .S1(_3131_),
    .X(_3500_));
 sky130_fd_sc_hd__mux2_1 _4396_ (.A0(_3066_),
    .A1(_3500_),
    .S(_3077_),
    .X(_3501_));
 sky130_fd_sc_hd__nor2_1 _4397_ (.A(_3108_),
    .B(_3501_),
    .Y(_3502_));
 sky130_fd_sc_hd__a211o_1 _4398_ (.A1(_3108_),
    .A2(_3056_),
    .B1(_3200_),
    .C1(_3502_),
    .X(_3503_));
 sky130_fd_sc_hd__o21ba_1 _4399_ (.A1(_1209_),
    .A2(_3480_),
    .B1_N(_3204_),
    .X(_3504_));
 sky130_fd_sc_hd__o22a_1 _4400_ (.A1(_0860_),
    .A2(_3503_),
    .B1(_3504_),
    .B2(_3481_),
    .X(_3505_));
 sky130_fd_sc_hd__or4b_1 _4401_ (.A(_3489_),
    .B(_3495_),
    .C(_3499_),
    .D_N(_3505_),
    .X(_3506_));
 sky130_fd_sc_hd__a31o_1 _4402_ (.A1(_2980_),
    .A2(_3484_),
    .A3(_3485_),
    .B1(_3506_),
    .X(_3507_));
 sky130_fd_sc_hd__a31o_2 _4403_ (.A1(_3305_),
    .A2(_3478_),
    .A3(_3479_),
    .B1(_3507_),
    .X(net100));
 sky130_fd_sc_hd__and3_1 _4404_ (.A(_1384_),
    .B(_3425_),
    .C(_3421_),
    .X(_3508_));
 sky130_fd_sc_hd__and2b_1 _4405_ (.A_N(_3437_),
    .B(_3429_),
    .X(_3509_));
 sky130_fd_sc_hd__and2_1 _4406_ (.A(_3428_),
    .B(_3438_),
    .X(_3510_));
 sky130_fd_sc_hd__clkbuf_4 _4407_ (.A(net34),
    .X(_3511_));
 sky130_fd_sc_hd__clkbuf_4 _4408_ (.A(_3511_),
    .X(_3512_));
 sky130_fd_sc_hd__clkbuf_4 _4409_ (.A(_3512_),
    .X(_3513_));
 sky130_fd_sc_hd__a22oi_1 _4410_ (.A1(_0445_),
    .A2(_3424_),
    .B1(_3513_),
    .B2(_0991_),
    .Y(_3514_));
 sky130_fd_sc_hd__and4_2 _4411_ (.A(_0707_),
    .B(_0477_),
    .C(_3424_),
    .D(_3512_),
    .X(_3515_));
 sky130_fd_sc_hd__nor2_1 _4412_ (.A(_3514_),
    .B(_3515_),
    .Y(_3516_));
 sky130_fd_sc_hd__o21ai_4 _4413_ (.A1(_3509_),
    .A2(_3510_),
    .B1(_3516_),
    .Y(_3517_));
 sky130_fd_sc_hd__or3_1 _4414_ (.A(_3509_),
    .B(_3510_),
    .C(_3516_),
    .X(_3518_));
 sky130_fd_sc_hd__and2_1 _4415_ (.A(_3517_),
    .B(_3518_),
    .X(_3519_));
 sky130_fd_sc_hd__and4_1 _4416_ (.A(_0205_),
    .B(_0335_),
    .C(_3196_),
    .D(_3272_),
    .X(_3520_));
 sky130_fd_sc_hd__nor2_1 _4417_ (.A(_3520_),
    .B(_3436_),
    .Y(_3521_));
 sky130_fd_sc_hd__o2bb2a_1 _4418_ (.A1_N(_2379_),
    .A2_N(_3443_),
    .B1(_3445_),
    .B2(_3441_),
    .X(_3522_));
 sky130_fd_sc_hd__a22o_1 _4419_ (.A1(_0085_),
    .A2(_3433_),
    .B1(_3431_),
    .B2(_1264_),
    .X(_3523_));
 sky130_fd_sc_hd__nand4_1 _4420_ (.A(_0085_),
    .B(_1264_),
    .C(_3195_),
    .D(_3431_),
    .Y(_3524_));
 sky130_fd_sc_hd__a22oi_1 _4421_ (.A1(_0739_),
    .A2(_3430_),
    .B1(_3523_),
    .B2(_3524_),
    .Y(_3525_));
 sky130_fd_sc_hd__and4_1 _4422_ (.A(_0324_),
    .B(_3343_),
    .C(_3523_),
    .D(_3524_),
    .X(_3526_));
 sky130_fd_sc_hd__or2_2 _4423_ (.A(_3525_),
    .B(_3526_),
    .X(_3527_));
 sky130_fd_sc_hd__xor2_1 _4424_ (.A(_3522_),
    .B(_3527_),
    .X(_3528_));
 sky130_fd_sc_hd__xnor2_1 _4425_ (.A(_3521_),
    .B(_3528_),
    .Y(_3529_));
 sky130_fd_sc_hd__buf_4 _4426_ (.A(_2423_),
    .X(_3530_));
 sky130_fd_sc_hd__clkbuf_4 _4427_ (.A(net59),
    .X(_3531_));
 sky130_fd_sc_hd__and3_1 _4428_ (.A(_0161_),
    .B(_3531_),
    .C(_2368_),
    .X(_3532_));
 sky130_fd_sc_hd__a22o_1 _4429_ (.A1(_3531_),
    .A2(_2368_),
    .B1(_2423_),
    .B2(_0161_),
    .X(_3533_));
 sky130_fd_sc_hd__a21bo_1 _4430_ (.A1(_3530_),
    .A2(_3532_),
    .B1_N(_3533_),
    .X(_3534_));
 sky130_fd_sc_hd__xnor2_2 _4431_ (.A(_2925_),
    .B(_3534_),
    .Y(_3535_));
 sky130_fd_sc_hd__and2_1 _4432_ (.A(_0292_),
    .B(_2106_),
    .X(_3536_));
 sky130_fd_sc_hd__clkbuf_4 _4433_ (.A(net2),
    .X(_3537_));
 sky130_fd_sc_hd__a22o_1 _4434_ (.A1(_3448_),
    .A2(net32),
    .B1(_3537_),
    .B2(_3449_),
    .X(_3538_));
 sky130_fd_sc_hd__nand4_2 _4435_ (.A(_3451_),
    .B(_3452_),
    .C(_2149_),
    .D(_2204_),
    .Y(_3539_));
 sky130_fd_sc_hd__nand3_1 _4436_ (.A(_3536_),
    .B(_3538_),
    .C(_3539_),
    .Y(_3540_));
 sky130_fd_sc_hd__a21o_1 _4437_ (.A1(_3538_),
    .A2(_3539_),
    .B1(_3536_),
    .X(_3541_));
 sky130_fd_sc_hd__a21bo_1 _4438_ (.A1(_3447_),
    .A2(_3450_),
    .B1_N(_3453_),
    .X(_3542_));
 sky130_fd_sc_hd__nand3_2 _4439_ (.A(_3540_),
    .B(_3541_),
    .C(_3542_),
    .Y(_3543_));
 sky130_fd_sc_hd__a21o_1 _4440_ (.A1(_3540_),
    .A2(_3541_),
    .B1(_3542_),
    .X(_3544_));
 sky130_fd_sc_hd__nand3_2 _4441_ (.A(_3535_),
    .B(_3543_),
    .C(_3544_),
    .Y(_3545_));
 sky130_fd_sc_hd__a21o_1 _4442_ (.A1(_3543_),
    .A2(_3544_),
    .B1(_3535_),
    .X(_3546_));
 sky130_fd_sc_hd__a21bo_1 _4443_ (.A1(_3446_),
    .A2(_3458_),
    .B1_N(_3457_),
    .X(_3547_));
 sky130_fd_sc_hd__nand3_2 _4444_ (.A(_3545_),
    .B(_3546_),
    .C(_3547_),
    .Y(_3548_));
 sky130_fd_sc_hd__a21o_1 _4445_ (.A1(_3545_),
    .A2(_3546_),
    .B1(_3547_),
    .X(_3549_));
 sky130_fd_sc_hd__and3_1 _4446_ (.A(net131),
    .B(_3548_),
    .C(_3549_),
    .X(_3550_));
 sky130_fd_sc_hd__a21oi_2 _4447_ (.A1(_3548_),
    .A2(_3549_),
    .B1(net131),
    .Y(_3551_));
 sky130_fd_sc_hd__a211o_2 _4448_ (.A1(_3462_),
    .A2(_3464_),
    .B1(_3550_),
    .C1(_3551_),
    .X(_3552_));
 sky130_fd_sc_hd__o211ai_4 _4449_ (.A1(_3550_),
    .A2(_3551_),
    .B1(_3462_),
    .C1(_3464_),
    .Y(_3553_));
 sky130_fd_sc_hd__and3_1 _4450_ (.A(_3519_),
    .B(_3552_),
    .C(_3553_),
    .X(_3554_));
 sky130_fd_sc_hd__a21oi_2 _4451_ (.A1(_3552_),
    .A2(_3553_),
    .B1(_3519_),
    .Y(_3555_));
 sky130_fd_sc_hd__a211o_1 _4452_ (.A1(_3466_),
    .A2(_3468_),
    .B1(_3554_),
    .C1(_3555_),
    .X(_3556_));
 sky130_fd_sc_hd__o211ai_4 _4453_ (.A1(_3554_),
    .A2(_3555_),
    .B1(_3466_),
    .C1(_3468_),
    .Y(_3557_));
 sky130_fd_sc_hd__and3_1 _4454_ (.A(_3508_),
    .B(_3556_),
    .C(_3557_),
    .X(_3558_));
 sky130_fd_sc_hd__a21oi_2 _4455_ (.A1(net144),
    .A2(_3557_),
    .B1(_3508_),
    .Y(_3559_));
 sky130_fd_sc_hd__a21o_1 _4456_ (.A1(_3377_),
    .A2(_3471_),
    .B1(_3470_),
    .X(_3560_));
 sky130_fd_sc_hd__or3_1 _4457_ (.A(_3558_),
    .B(_3559_),
    .C(_3560_),
    .X(_3561_));
 sky130_fd_sc_hd__o21ai_2 _4458_ (.A1(_3558_),
    .A2(_3559_),
    .B1(_3560_),
    .Y(_3562_));
 sky130_fd_sc_hd__or2_1 _4459_ (.A(_3379_),
    .B(_3472_),
    .X(_3563_));
 sky130_fd_sc_hd__a21o_1 _4460_ (.A1(_3561_),
    .A2(_3562_),
    .B1(_3563_),
    .X(_3564_));
 sky130_fd_sc_hd__nand3_1 _4461_ (.A(_3563_),
    .B(_3561_),
    .C(_3562_),
    .Y(_3565_));
 sky130_fd_sc_hd__and3_1 _4462_ (.A(_3476_),
    .B(_3564_),
    .C(_3565_),
    .X(_3566_));
 sky130_fd_sc_hd__a21oi_1 _4463_ (.A1(_3564_),
    .A2(_3565_),
    .B1(_3476_),
    .Y(_3567_));
 sky130_fd_sc_hd__or2_1 _4464_ (.A(_3566_),
    .B(_3567_),
    .X(_3568_));
 sky130_fd_sc_hd__nand2_1 _4465_ (.A(_3479_),
    .B(_3568_),
    .Y(_3569_));
 sky130_fd_sc_hd__o21a_1 _4466_ (.A1(_3479_),
    .A2(_3568_),
    .B1(_3305_),
    .X(_3570_));
 sky130_fd_sc_hd__buf_4 _4467_ (.A(_0652_),
    .X(_3571_));
 sky130_fd_sc_hd__buf_2 _4468_ (.A(net34),
    .X(_3572_));
 sky130_fd_sc_hd__and2_4 _4469_ (.A(net2),
    .B(_3572_),
    .X(_3573_));
 sky130_fd_sc_hd__nor2_1 _4470_ (.A(_2237_),
    .B(_3513_),
    .Y(_3574_));
 sky130_fd_sc_hd__or2_2 _4471_ (.A(_3573_),
    .B(_3574_),
    .X(_3575_));
 sky130_fd_sc_hd__and2b_1 _4472_ (.A_N(_3425_),
    .B(_2182_),
    .X(_3576_));
 sky130_fd_sc_hd__a21o_1 _4473_ (.A1(_3482_),
    .A2(_3497_),
    .B1(_3576_),
    .X(_3577_));
 sky130_fd_sc_hd__or2_1 _4474_ (.A(_3575_),
    .B(_3577_),
    .X(_3578_));
 sky130_fd_sc_hd__nand2_1 _4475_ (.A(_3575_),
    .B(_3577_),
    .Y(_3579_));
 sky130_fd_sc_hd__buf_2 _4476_ (.A(_3127_),
    .X(_3580_));
 sky130_fd_sc_hd__mux2_1 _4477_ (.A0(_3220_),
    .A1(_3221_),
    .S(_3077_),
    .X(_3581_));
 sky130_fd_sc_hd__mux2_1 _4478_ (.A0(_3219_),
    .A1(_3225_),
    .S(_1100_),
    .X(_3582_));
 sky130_fd_sc_hd__mux2_1 _4479_ (.A0(_3581_),
    .A1(_3582_),
    .S(_3486_),
    .X(_3583_));
 sky130_fd_sc_hd__a22o_1 _4480_ (.A1(_2062_),
    .A2(_3024_),
    .B1(_3224_),
    .B2(_3077_),
    .X(_3584_));
 sky130_fd_sc_hd__nand2_1 _4481_ (.A(_3301_),
    .B(_3584_),
    .Y(_3585_));
 sky130_fd_sc_hd__nand2_1 _4482_ (.A(_3580_),
    .B(_3585_),
    .Y(_3586_));
 sky130_fd_sc_hd__clkbuf_4 _4483_ (.A(_1701_),
    .X(_3587_));
 sky130_fd_sc_hd__o211a_1 _4484_ (.A1(_3580_),
    .A2(_3583_),
    .B1(_3586_),
    .C1(_3587_),
    .X(_3588_));
 sky130_fd_sc_hd__clkbuf_4 _4485_ (.A(_1209_),
    .X(_3589_));
 sky130_fd_sc_hd__o21ba_1 _4486_ (.A1(_3589_),
    .A2(_3573_),
    .B1_N(_3204_),
    .X(_3590_));
 sky130_fd_sc_hd__clkbuf_4 _4487_ (.A(_0969_),
    .X(_3591_));
 sky130_fd_sc_hd__a21o_1 _4488_ (.A1(_3490_),
    .A2(_3591_),
    .B1(_3486_),
    .X(_3592_));
 sky130_fd_sc_hd__a2bb2o_1 _4489_ (.A1_N(_3574_),
    .A2_N(_3590_),
    .B1(_3592_),
    .B2(_3201_),
    .X(_3593_));
 sky130_fd_sc_hd__a221o_1 _4490_ (.A1(_3194_),
    .A2(_3573_),
    .B1(_3574_),
    .B2(_3414_),
    .C1(_3593_),
    .X(_3594_));
 sky130_fd_sc_hd__or2_1 _4491_ (.A(_0783_),
    .B(_0641_),
    .X(_3595_));
 sky130_fd_sc_hd__clkbuf_4 _4492_ (.A(_3595_),
    .X(_3596_));
 sky130_fd_sc_hd__o211a_1 _4493_ (.A1(_2182_),
    .A2(_3425_),
    .B1(_2138_),
    .C1(_3386_),
    .X(_3597_));
 sky130_fd_sc_hd__nor2_1 _4494_ (.A(_3480_),
    .B(_3597_),
    .Y(_3598_));
 sky130_fd_sc_hd__a211o_1 _4495_ (.A1(_3395_),
    .A2(_3396_),
    .B1(_3482_),
    .C1(_3389_),
    .X(_3599_));
 sky130_fd_sc_hd__and3_1 _4496_ (.A(_3575_),
    .B(_3598_),
    .C(_3599_),
    .X(_3600_));
 sky130_fd_sc_hd__a21oi_2 _4497_ (.A1(_3598_),
    .A2(_3599_),
    .B1(_3575_),
    .Y(_3601_));
 sky130_fd_sc_hd__mux4_1 _4498_ (.A0(_2237_),
    .A1(_2182_),
    .A2(_2138_),
    .A3(_3139_),
    .S0(_0925_),
    .S1(_0969_),
    .X(_3602_));
 sky130_fd_sc_hd__mux2_1 _4499_ (.A0(_3207_),
    .A1(_3602_),
    .S(_3077_),
    .X(_3603_));
 sky130_fd_sc_hd__mux2_1 _4500_ (.A0(_3212_),
    .A1(_3603_),
    .S(_3301_),
    .X(_3604_));
 sky130_fd_sc_hd__or2b_1 _4501_ (.A(_1734_),
    .B_N(_3604_),
    .X(_3605_));
 sky130_fd_sc_hd__o32a_1 _4502_ (.A1(_3596_),
    .A2(_3600_),
    .A3(_3601_),
    .B1(_3605_),
    .B2(_0860_),
    .X(_3606_));
 sky130_fd_sc_hd__or3b_1 _4503_ (.A(_3588_),
    .B(_3594_),
    .C_N(_3606_),
    .X(_3607_));
 sky130_fd_sc_hd__a31o_1 _4504_ (.A1(_3571_),
    .A2(_3578_),
    .A3(_3579_),
    .B1(_3607_),
    .X(_3608_));
 sky130_fd_sc_hd__a21o_2 _4505_ (.A1(_3569_),
    .A2(_3570_),
    .B1(_3608_),
    .X(net70));
 sky130_fd_sc_hd__a21oi_1 _4506_ (.A1(_3561_),
    .A2(_3562_),
    .B1(_3563_),
    .Y(_3609_));
 sky130_fd_sc_hd__o21ba_1 _4507_ (.A1(_3479_),
    .A2(_3567_),
    .B1_N(_3566_),
    .X(_3610_));
 sky130_fd_sc_hd__nand3_2 _4508_ (.A(_3508_),
    .B(net144),
    .C(_3557_),
    .Y(_3611_));
 sky130_fd_sc_hd__and3b_1 _4509_ (.A_N(_3559_),
    .B(_3470_),
    .C(_3611_),
    .X(_3612_));
 sky130_fd_sc_hd__nand3_2 _4510_ (.A(_3519_),
    .B(_3552_),
    .C(_3553_),
    .Y(_3613_));
 sky130_fd_sc_hd__or2b_1 _4511_ (.A(_3521_),
    .B_N(_3528_),
    .X(_3614_));
 sky130_fd_sc_hd__o21ai_2 _4512_ (.A1(_3522_),
    .A2(_3527_),
    .B1(_3614_),
    .Y(_3615_));
 sky130_fd_sc_hd__and4_1 _4513_ (.A(_0314_),
    .B(_0412_),
    .C(net64),
    .D(_3572_),
    .X(_3616_));
 sky130_fd_sc_hd__a22o_1 _4514_ (.A1(_0314_),
    .A2(net64),
    .B1(_3572_),
    .B2(net163),
    .X(_3617_));
 sky130_fd_sc_hd__and4b_1 _4515_ (.A_N(_3616_),
    .B(net35),
    .C(net1),
    .D(_3617_),
    .X(_3618_));
 sky130_fd_sc_hd__buf_2 _4516_ (.A(net35),
    .X(_3619_));
 sky130_fd_sc_hd__buf_4 _4517_ (.A(_3619_),
    .X(_3620_));
 sky130_fd_sc_hd__inv_2 _4518_ (.A(_3616_),
    .Y(_3621_));
 sky130_fd_sc_hd__a22oi_1 _4519_ (.A1(_0477_),
    .A2(_3620_),
    .B1(_3617_),
    .B2(_3621_),
    .Y(_3622_));
 sky130_fd_sc_hd__nor2_1 _4520_ (.A(_3618_),
    .B(_3622_),
    .Y(_3623_));
 sky130_fd_sc_hd__and2_1 _4521_ (.A(_3515_),
    .B(_3623_),
    .X(_3624_));
 sky130_fd_sc_hd__nor2_1 _4522_ (.A(_3515_),
    .B(_3623_),
    .Y(_3625_));
 sky130_fd_sc_hd__or2_1 _4523_ (.A(_3624_),
    .B(_3625_),
    .X(_3626_));
 sky130_fd_sc_hd__xnor2_1 _4524_ (.A(_3615_),
    .B(_3626_),
    .Y(_3627_));
 sky130_fd_sc_hd__nand3_1 _4525_ (.A(_3529_),
    .B(_3548_),
    .C(_3549_),
    .Y(_3628_));
 sky130_fd_sc_hd__a41o_2 _4526_ (.A1(_0106_),
    .A2(_0215_),
    .A3(_3197_),
    .A4(_3272_),
    .B1(_3526_),
    .X(_3629_));
 sky130_fd_sc_hd__a22o_1 _4527_ (.A1(_2925_),
    .A2(_3533_),
    .B1(_3532_),
    .B2(_3530_),
    .X(_3630_));
 sky130_fd_sc_hd__clkbuf_4 _4528_ (.A(_3343_),
    .X(_3631_));
 sky130_fd_sc_hd__buf_4 _4529_ (.A(net61),
    .X(_3632_));
 sky130_fd_sc_hd__clkbuf_4 _4530_ (.A(_3270_),
    .X(_3633_));
 sky130_fd_sc_hd__a22o_1 _4531_ (.A1(_2302_),
    .A2(_3632_),
    .B1(_3633_),
    .B2(_0085_),
    .X(_3634_));
 sky130_fd_sc_hd__clkbuf_4 _4532_ (.A(net28),
    .X(_3635_));
 sky130_fd_sc_hd__nand4_2 _4533_ (.A(_3440_),
    .B(_3635_),
    .C(_3632_),
    .D(_3271_),
    .Y(_3636_));
 sky130_fd_sc_hd__nand4_2 _4534_ (.A(_0205_),
    .B(_3631_),
    .C(_3634_),
    .D(_3636_),
    .Y(_3637_));
 sky130_fd_sc_hd__a22o_1 _4535_ (.A1(_1275_),
    .A2(_3631_),
    .B1(_3634_),
    .B2(_3636_),
    .X(_3638_));
 sky130_fd_sc_hd__and3_1 _4536_ (.A(_3630_),
    .B(_3637_),
    .C(_3638_),
    .X(_3639_));
 sky130_fd_sc_hd__a21oi_1 _4537_ (.A1(_3637_),
    .A2(_3638_),
    .B1(_3630_),
    .Y(_3640_));
 sky130_fd_sc_hd__nor2_1 _4538_ (.A(_3639_),
    .B(_3640_),
    .Y(_3641_));
 sky130_fd_sc_hd__xor2_2 _4539_ (.A(_3629_),
    .B(_3641_),
    .X(_3642_));
 sky130_fd_sc_hd__nand2_1 _4540_ (.A(_2881_),
    .B(_2379_),
    .Y(_3643_));
 sky130_fd_sc_hd__buf_4 _4541_ (.A(net31),
    .X(_3644_));
 sky130_fd_sc_hd__buf_4 _4542_ (.A(_3169_),
    .X(_3645_));
 sky130_fd_sc_hd__a22oi_2 _4543_ (.A1(_0041_),
    .A2(_2434_),
    .B1(_3644_),
    .B2(_3645_),
    .Y(_3646_));
 sky130_fd_sc_hd__and4_1 _4544_ (.A(_3645_),
    .B(_3531_),
    .C(_2434_),
    .D(_2106_),
    .X(_3647_));
 sky130_fd_sc_hd__nor2_1 _4545_ (.A(_3646_),
    .B(_3647_),
    .Y(_3648_));
 sky130_fd_sc_hd__xnor2_1 _4546_ (.A(_3643_),
    .B(_3648_),
    .Y(_3649_));
 sky130_fd_sc_hd__and2_1 _4547_ (.A(_0292_),
    .B(net32),
    .X(_3650_));
 sky130_fd_sc_hd__clkbuf_4 _4548_ (.A(net3),
    .X(_3651_));
 sky130_fd_sc_hd__a22o_1 _4549_ (.A1(_3448_),
    .A2(_3537_),
    .B1(_3651_),
    .B2(_3449_),
    .X(_3652_));
 sky130_fd_sc_hd__nand4_2 _4550_ (.A(_3451_),
    .B(_3452_),
    .C(_3537_),
    .D(_3651_),
    .Y(_3653_));
 sky130_fd_sc_hd__nand3_1 _4551_ (.A(_3650_),
    .B(_3652_),
    .C(_3653_),
    .Y(_3654_));
 sky130_fd_sc_hd__a21o_1 _4552_ (.A1(_3652_),
    .A2(_3653_),
    .B1(_3650_),
    .X(_3655_));
 sky130_fd_sc_hd__a21bo_1 _4553_ (.A1(_3536_),
    .A2(_3538_),
    .B1_N(_3539_),
    .X(_3656_));
 sky130_fd_sc_hd__nand3_1 _4554_ (.A(_3654_),
    .B(_3655_),
    .C(_3656_),
    .Y(_3657_));
 sky130_fd_sc_hd__a21o_1 _4555_ (.A1(_3654_),
    .A2(_3655_),
    .B1(_3656_),
    .X(_3658_));
 sky130_fd_sc_hd__nand3_1 _4556_ (.A(_3649_),
    .B(_3657_),
    .C(_3658_),
    .Y(_3659_));
 sky130_fd_sc_hd__a21o_1 _4557_ (.A1(_3657_),
    .A2(_3658_),
    .B1(_3649_),
    .X(_3660_));
 sky130_fd_sc_hd__a21bo_1 _4558_ (.A1(_3535_),
    .A2(_3544_),
    .B1_N(_3543_),
    .X(_3661_));
 sky130_fd_sc_hd__nand3_2 _4559_ (.A(_3659_),
    .B(_3660_),
    .C(_3661_),
    .Y(_3662_));
 sky130_fd_sc_hd__a21o_1 _4560_ (.A1(_3659_),
    .A2(_3660_),
    .B1(_3661_),
    .X(_3663_));
 sky130_fd_sc_hd__and3_1 _4561_ (.A(_3642_),
    .B(_3662_),
    .C(_3663_),
    .X(_3664_));
 sky130_fd_sc_hd__a21oi_2 _4562_ (.A1(_3662_),
    .A2(_3663_),
    .B1(_3642_),
    .Y(_3665_));
 sky130_fd_sc_hd__a211o_1 _4563_ (.A1(_3548_),
    .A2(_3628_),
    .B1(_3664_),
    .C1(_3665_),
    .X(_3666_));
 sky130_fd_sc_hd__o211ai_2 _4564_ (.A1(_3664_),
    .A2(_3665_),
    .B1(_3548_),
    .C1(net155),
    .Y(_3667_));
 sky130_fd_sc_hd__and3_2 _4565_ (.A(_3627_),
    .B(_3666_),
    .C(_3667_),
    .X(_3668_));
 sky130_fd_sc_hd__a21oi_2 _4566_ (.A1(net139),
    .A2(_3667_),
    .B1(_3627_),
    .Y(_3669_));
 sky130_fd_sc_hd__a211oi_4 _4567_ (.A1(_3552_),
    .A2(_3613_),
    .B1(_3668_),
    .C1(_3669_),
    .Y(_3670_));
 sky130_fd_sc_hd__o211a_1 _4568_ (.A1(_3668_),
    .A2(_3669_),
    .B1(_3552_),
    .C1(_3613_),
    .X(_3671_));
 sky130_fd_sc_hd__nor3_4 _4569_ (.A(_3517_),
    .B(_3670_),
    .C(_3671_),
    .Y(_3672_));
 sky130_fd_sc_hd__o21a_1 _4570_ (.A1(_3670_),
    .A2(_3671_),
    .B1(_3517_),
    .X(_3673_));
 sky130_fd_sc_hd__a211o_1 _4571_ (.A1(net144),
    .A2(_3611_),
    .B1(_3672_),
    .C1(_3673_),
    .X(_3674_));
 sky130_fd_sc_hd__o211ai_4 _4572_ (.A1(_3672_),
    .A2(_3673_),
    .B1(net144),
    .C1(_3611_),
    .Y(_3675_));
 sky130_fd_sc_hd__and3_1 _4573_ (.A(_3612_),
    .B(_3674_),
    .C(_3675_),
    .X(_3676_));
 sky130_fd_sc_hd__a21oi_1 _4574_ (.A1(_3674_),
    .A2(_3675_),
    .B1(_3612_),
    .Y(_3677_));
 sky130_fd_sc_hd__or4_1 _4575_ (.A(_3473_),
    .B(_3472_),
    .C(_3558_),
    .D(_3559_),
    .X(_3678_));
 sky130_fd_sc_hd__or3_1 _4576_ (.A(_3676_),
    .B(_3677_),
    .C(_3678_),
    .X(_3679_));
 sky130_fd_sc_hd__o21ai_1 _4577_ (.A1(_3676_),
    .A2(_3677_),
    .B1(_3678_),
    .Y(_3680_));
 sky130_fd_sc_hd__nand2_1 _4578_ (.A(_3679_),
    .B(_3680_),
    .Y(_3681_));
 sky130_fd_sc_hd__xor2_1 _4579_ (.A(_3610_),
    .B(_3681_),
    .X(_3682_));
 sky130_fd_sc_hd__or2_1 _4580_ (.A(_3609_),
    .B(net126),
    .X(_3683_));
 sky130_fd_sc_hd__nand2_1 _4581_ (.A(_3609_),
    .B(net127),
    .Y(_3684_));
 sky130_fd_sc_hd__clkbuf_4 _4582_ (.A(_3620_),
    .X(_3685_));
 sky130_fd_sc_hd__or2_1 _4583_ (.A(_2270_),
    .B(_3685_),
    .X(_3686_));
 sky130_fd_sc_hd__nand2_1 _4584_ (.A(_3137_),
    .B(_3685_),
    .Y(_3687_));
 sky130_fd_sc_hd__nand2_1 _4585_ (.A(_3686_),
    .B(_3687_),
    .Y(_3688_));
 sky130_fd_sc_hd__and2b_1 _4586_ (.A_N(_3513_),
    .B(_2237_),
    .X(_3689_));
 sky130_fd_sc_hd__a21o_1 _4587_ (.A1(_3575_),
    .A2(_3577_),
    .B1(_3689_),
    .X(_3690_));
 sky130_fd_sc_hd__or2_1 _4588_ (.A(_3688_),
    .B(_3690_),
    .X(_3691_));
 sky130_fd_sc_hd__and2_1 _4589_ (.A(_3688_),
    .B(_3690_),
    .X(_3692_));
 sky130_fd_sc_hd__inv_2 _4590_ (.A(_3692_),
    .Y(_3693_));
 sky130_fd_sc_hd__or3b_1 _4591_ (.A(_3573_),
    .B(_3601_),
    .C_N(_3688_),
    .X(_3694_));
 sky130_fd_sc_hd__o21ba_1 _4592_ (.A1(_3573_),
    .A2(_3601_),
    .B1_N(_3688_),
    .X(_3695_));
 sky130_fd_sc_hd__inv_2 _4593_ (.A(_3695_),
    .Y(_3696_));
 sky130_fd_sc_hd__mux4_1 _4594_ (.A0(_3296_),
    .A1(_3299_),
    .A2(_3292_),
    .A3(_3298_),
    .S0(_3301_),
    .S1(_3490_),
    .X(_3697_));
 sky130_fd_sc_hd__o2bb2a_1 _4595_ (.A1_N(_0554_),
    .A2_N(_3291_),
    .B1(_3035_),
    .B2(_3144_),
    .X(_3698_));
 sky130_fd_sc_hd__or2_2 _4596_ (.A(_3108_),
    .B(_3698_),
    .X(_3699_));
 sky130_fd_sc_hd__nand2_1 _4597_ (.A(_3127_),
    .B(_3699_),
    .Y(_3700_));
 sky130_fd_sc_hd__o211a_1 _4598_ (.A1(_3580_),
    .A2(_3697_),
    .B1(_3700_),
    .C1(_3587_),
    .X(_3701_));
 sky130_fd_sc_hd__mux4_1 _4599_ (.A0(_3137_),
    .A1(_2237_),
    .A2(_2182_),
    .A3(_2138_),
    .S0(_3046_),
    .S1(_3591_),
    .X(_3702_));
 sky130_fd_sc_hd__mux2_1 _4600_ (.A0(_3283_),
    .A1(_3702_),
    .S(_3087_),
    .X(_3703_));
 sky130_fd_sc_hd__a21o_1 _4601_ (.A1(_3087_),
    .A2(_3284_),
    .B1(_3301_),
    .X(_3704_));
 sky130_fd_sc_hd__o21ai_2 _4602_ (.A1(_3486_),
    .A2(_3703_),
    .B1(_3704_),
    .Y(_3705_));
 sky130_fd_sc_hd__nor2_1 _4603_ (.A(_0860_),
    .B(_3705_),
    .Y(_3706_));
 sky130_fd_sc_hd__o21a_1 _4604_ (.A1(_3046_),
    .A2(_3591_),
    .B1(_3490_),
    .X(_3707_));
 sky130_fd_sc_hd__o21a_1 _4605_ (.A1(_3486_),
    .A2(_3707_),
    .B1(_3201_),
    .X(_3708_));
 sky130_fd_sc_hd__and2_2 _4606_ (.A(_2248_),
    .B(net35),
    .X(_3709_));
 sky130_fd_sc_hd__a21o_1 _4607_ (.A1(net124),
    .A2(_3687_),
    .B1(_3204_),
    .X(_3710_));
 sky130_fd_sc_hd__or4b_1 _4608_ (.A(_1165_),
    .B(_0630_),
    .C(_1144_),
    .D_N(_1154_),
    .X(_3711_));
 sky130_fd_sc_hd__clkbuf_4 _4609_ (.A(_3711_),
    .X(_3712_));
 sky130_fd_sc_hd__nor2_1 _4610_ (.A(_3712_),
    .B(_3686_),
    .Y(_3713_));
 sky130_fd_sc_hd__a221o_1 _4611_ (.A1(_3194_),
    .A2(_3709_),
    .B1(_3710_),
    .B2(_3686_),
    .C1(_3713_),
    .X(_3714_));
 sky130_fd_sc_hd__or4_1 _4612_ (.A(_3701_),
    .B(_3706_),
    .C(_3708_),
    .D(_3714_),
    .X(_3715_));
 sky130_fd_sc_hd__a31o_1 _4613_ (.A1(_2980_),
    .A2(_3694_),
    .A3(_3696_),
    .B1(_3715_),
    .X(_3716_));
 sky130_fd_sc_hd__a31o_1 _4614_ (.A1(_0652_),
    .A2(_3691_),
    .A3(_3693_),
    .B1(_3716_),
    .X(_3717_));
 sky130_fd_sc_hd__a31o_2 _4615_ (.A1(_3305_),
    .A2(_3683_),
    .A3(_3684_),
    .B1(_3717_),
    .X(net71));
 sky130_fd_sc_hd__buf_2 _4616_ (.A(net36),
    .X(_3718_));
 sky130_fd_sc_hd__clkbuf_4 _4617_ (.A(_3718_),
    .X(_3719_));
 sky130_fd_sc_hd__clkbuf_4 _4618_ (.A(_3719_),
    .X(_3720_));
 sky130_fd_sc_hd__nor2_1 _4619_ (.A(_2675_),
    .B(_3720_),
    .Y(_3721_));
 sky130_fd_sc_hd__and2_2 _4620_ (.A(_2653_),
    .B(_3718_),
    .X(_3722_));
 sky130_fd_sc_hd__or2_1 _4621_ (.A(_3721_),
    .B(_3722_),
    .X(_3723_));
 sky130_fd_sc_hd__o21ba_1 _4622_ (.A1(_3709_),
    .A2(_3695_),
    .B1_N(_3723_),
    .X(_3724_));
 sky130_fd_sc_hd__or2_1 _4623_ (.A(_3596_),
    .B(_3724_),
    .X(_3725_));
 sky130_fd_sc_hd__a31oi_1 _4624_ (.A1(_3687_),
    .A2(_3696_),
    .A3(_3723_),
    .B1(_3725_),
    .Y(_3726_));
 sky130_fd_sc_hd__buf_2 _4625_ (.A(_3580_),
    .X(_3727_));
 sky130_fd_sc_hd__mux4_1 _4626_ (.A0(_1843_),
    .A1(_1985_),
    .A2(_2631_),
    .A3(_2806_),
    .S0(_3087_),
    .S1(_3301_),
    .X(_3728_));
 sky130_fd_sc_hd__nor2_1 _4627_ (.A(_0980_),
    .B(_0870_),
    .Y(_3729_));
 sky130_fd_sc_hd__nand2_1 _4628_ (.A(_2073_),
    .B(_3729_),
    .Y(_3730_));
 sky130_fd_sc_hd__nand2_1 _4629_ (.A(_3727_),
    .B(_3730_),
    .Y(_3731_));
 sky130_fd_sc_hd__o211a_1 _4630_ (.A1(_3727_),
    .A2(_3728_),
    .B1(_3731_),
    .C1(_3587_),
    .X(_3732_));
 sky130_fd_sc_hd__buf_2 _4631_ (.A(_3204_),
    .X(_0000_));
 sky130_fd_sc_hd__o21ba_1 _4632_ (.A1(_3589_),
    .A2(_3722_),
    .B1_N(_0000_),
    .X(_0001_));
 sky130_fd_sc_hd__or2_1 _4633_ (.A(_3490_),
    .B(_3486_),
    .X(_0002_));
 sky130_fd_sc_hd__inv_2 _4634_ (.A(_1111_),
    .Y(_0003_));
 sky130_fd_sc_hd__mux4_2 _4635_ (.A0(_2675_),
    .A1(_3137_),
    .A2(_2237_),
    .A3(_2182_),
    .S0(_3046_),
    .S1(_3591_),
    .X(_0004_));
 sky130_fd_sc_hd__mux2_1 _4636_ (.A0(_3407_),
    .A1(_0004_),
    .S(_3087_),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_1 _4637_ (.A0(_0003_),
    .A1(_0005_),
    .S(_3301_),
    .X(_0006_));
 sky130_fd_sc_hd__nor2_1 _4638_ (.A(_3580_),
    .B(_3118_),
    .Y(_0007_));
 sky130_fd_sc_hd__a22o_1 _4639_ (.A1(_3414_),
    .A2(_3721_),
    .B1(_3722_),
    .B2(_3194_),
    .X(_0008_));
 sky130_fd_sc_hd__a221o_1 _4640_ (.A1(_3201_),
    .A2(_0002_),
    .B1(_0006_),
    .B2(_0007_),
    .C1(_0008_),
    .X(_0009_));
 sky130_fd_sc_hd__o21bai_1 _4641_ (.A1(_3721_),
    .A2(_0001_),
    .B1_N(_0009_),
    .Y(_0010_));
 sky130_fd_sc_hd__and2b_1 _4642_ (.A_N(_3685_),
    .B(_3137_),
    .X(_0011_));
 sky130_fd_sc_hd__a21o_1 _4643_ (.A1(_3688_),
    .A2(_3690_),
    .B1(_0011_),
    .X(_0012_));
 sky130_fd_sc_hd__or2_1 _4644_ (.A(_3723_),
    .B(_0012_),
    .X(_0013_));
 sky130_fd_sc_hd__nand2_1 _4645_ (.A(_3723_),
    .B(_0012_),
    .Y(_0014_));
 sky130_fd_sc_hd__and2b_1 _4646_ (.A_N(_3626_),
    .B(_3615_),
    .X(_0015_));
 sky130_fd_sc_hd__inv_2 _4647_ (.A(_0015_),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _4648_ (.A(net138),
    .Y(_0017_));
 sky130_fd_sc_hd__a21oi_2 _4649_ (.A1(_3629_),
    .A2(_3641_),
    .B1(_3639_),
    .Y(_0018_));
 sky130_fd_sc_hd__nand2_1 _4650_ (.A(_0477_),
    .B(_3719_),
    .Y(_0019_));
 sky130_fd_sc_hd__a22oi_1 _4651_ (.A1(_0194_),
    .A2(_3422_),
    .B1(_3511_),
    .B2(_0324_),
    .Y(_0020_));
 sky130_fd_sc_hd__and4_1 _4652_ (.A(_1264_),
    .B(_0314_),
    .C(net64),
    .D(_3572_),
    .X(_0021_));
 sky130_fd_sc_hd__and4bb_1 _4653_ (.A_N(_0020_),
    .B_N(_0021_),
    .C(_0423_),
    .D(net35),
    .X(_0022_));
 sky130_fd_sc_hd__o2bb2a_1 _4654_ (.A1_N(_0423_),
    .A2_N(_3619_),
    .B1(_0020_),
    .B2(_0021_),
    .X(_0023_));
 sky130_fd_sc_hd__nor2_1 _4655_ (.A(_0022_),
    .B(_0023_),
    .Y(_0024_));
 sky130_fd_sc_hd__or2_1 _4656_ (.A(_3616_),
    .B(_3618_),
    .X(_0025_));
 sky130_fd_sc_hd__xor2_1 _4657_ (.A(_0024_),
    .B(_0025_),
    .X(_0026_));
 sky130_fd_sc_hd__xnor2_1 _4658_ (.A(_0019_),
    .B(_0026_),
    .Y(_0027_));
 sky130_fd_sc_hd__xnor2_1 _4659_ (.A(_0018_),
    .B(_0027_),
    .Y(_0028_));
 sky130_fd_sc_hd__xnor2_1 _4660_ (.A(_3624_),
    .B(_0028_),
    .Y(_0029_));
 sky130_fd_sc_hd__nand3_1 _4661_ (.A(_3642_),
    .B(_3662_),
    .C(_3663_),
    .Y(_0031_));
 sky130_fd_sc_hd__nand2_2 _4662_ (.A(_3636_),
    .B(_3637_),
    .Y(_0032_));
 sky130_fd_sc_hd__o21ba_1 _4663_ (.A1(_3643_),
    .A2(_3646_),
    .B1_N(_3647_),
    .X(_0033_));
 sky130_fd_sc_hd__nand2_1 _4664_ (.A(_0095_),
    .B(_3631_),
    .Y(_0034_));
 sky130_fd_sc_hd__and3_1 _4665_ (.A(_2368_),
    .B(_3433_),
    .C(_3431_),
    .X(_0035_));
 sky130_fd_sc_hd__a22o_1 _4666_ (.A1(_2368_),
    .A2(_3433_),
    .B1(_3431_),
    .B2(_2302_),
    .X(_0036_));
 sky130_fd_sc_hd__a21bo_1 _4667_ (.A1(_3635_),
    .A2(_0035_),
    .B1_N(_0036_),
    .X(_0037_));
 sky130_fd_sc_hd__xor2_2 _4668_ (.A(_0034_),
    .B(_0037_),
    .X(_0038_));
 sky130_fd_sc_hd__xnor2_2 _4669_ (.A(_0033_),
    .B(_0038_),
    .Y(_0039_));
 sky130_fd_sc_hd__xor2_2 _4670_ (.A(_0032_),
    .B(_0039_),
    .X(_0040_));
 sky130_fd_sc_hd__clkbuf_4 _4671_ (.A(net60),
    .X(_0042_));
 sky130_fd_sc_hd__nand2_1 _4672_ (.A(_0042_),
    .B(_3530_),
    .Y(_0043_));
 sky130_fd_sc_hd__a22oi_2 _4673_ (.A1(_0041_),
    .A2(_2106_),
    .B1(_2149_),
    .B2(_3645_),
    .Y(_0044_));
 sky130_fd_sc_hd__and4_1 _4674_ (.A(_0161_),
    .B(_3531_),
    .C(_2106_),
    .D(net32),
    .X(_0045_));
 sky130_fd_sc_hd__nor2_1 _4675_ (.A(_0044_),
    .B(_0045_),
    .Y(_0046_));
 sky130_fd_sc_hd__xnor2_2 _4676_ (.A(_0043_),
    .B(_0046_),
    .Y(_0047_));
 sky130_fd_sc_hd__and2_1 _4677_ (.A(_0281_),
    .B(_3537_),
    .X(_0048_));
 sky130_fd_sc_hd__a22o_1 _4678_ (.A1(_0390_),
    .A2(_3651_),
    .B1(_2642_),
    .B2(_0488_),
    .X(_0049_));
 sky130_fd_sc_hd__nand4_1 _4679_ (.A(_3449_),
    .B(_3448_),
    .C(_3651_),
    .D(_2642_),
    .Y(_0050_));
 sky130_fd_sc_hd__nand3_1 _4680_ (.A(_0048_),
    .B(_0049_),
    .C(_0050_),
    .Y(_0051_));
 sky130_fd_sc_hd__a21o_1 _4681_ (.A1(_0049_),
    .A2(_0050_),
    .B1(_0048_),
    .X(_0053_));
 sky130_fd_sc_hd__a21bo_1 _4682_ (.A1(_3650_),
    .A2(_3652_),
    .B1_N(_3653_),
    .X(_0054_));
 sky130_fd_sc_hd__nand3_1 _4683_ (.A(_0051_),
    .B(_0053_),
    .C(_0054_),
    .Y(_0055_));
 sky130_fd_sc_hd__a21o_1 _4684_ (.A1(_0051_),
    .A2(_0053_),
    .B1(_0054_),
    .X(_0056_));
 sky130_fd_sc_hd__nand3_2 _4685_ (.A(_0047_),
    .B(_0055_),
    .C(_0056_),
    .Y(_0057_));
 sky130_fd_sc_hd__a21o_1 _4686_ (.A1(_0055_),
    .A2(_0056_),
    .B1(_0047_),
    .X(_0058_));
 sky130_fd_sc_hd__a21bo_1 _4687_ (.A1(_3649_),
    .A2(_3658_),
    .B1_N(_3657_),
    .X(_0059_));
 sky130_fd_sc_hd__nand3_4 _4688_ (.A(_0057_),
    .B(_0058_),
    .C(_0059_),
    .Y(_0060_));
 sky130_fd_sc_hd__a21o_1 _4689_ (.A1(_0057_),
    .A2(_0058_),
    .B1(_0059_),
    .X(_0061_));
 sky130_fd_sc_hd__and3_1 _4690_ (.A(_0040_),
    .B(_0060_),
    .C(_0061_),
    .X(_0062_));
 sky130_fd_sc_hd__a21oi_1 _4691_ (.A1(_0060_),
    .A2(_0061_),
    .B1(_0040_),
    .Y(_0064_));
 sky130_fd_sc_hd__a211oi_2 _4692_ (.A1(_3662_),
    .A2(_0031_),
    .B1(_0062_),
    .C1(_0064_),
    .Y(_0065_));
 sky130_fd_sc_hd__o211a_1 _4693_ (.A1(_0062_),
    .A2(_0064_),
    .B1(_3662_),
    .C1(_0031_),
    .X(_0066_));
 sky130_fd_sc_hd__or3_2 _4694_ (.A(_0029_),
    .B(_0065_),
    .C(_0066_),
    .X(_0067_));
 sky130_fd_sc_hd__o21ai_1 _4695_ (.A1(_0065_),
    .A2(_0066_),
    .B1(_0029_),
    .Y(_0068_));
 sky130_fd_sc_hd__o211a_1 _4696_ (.A1(_0017_),
    .A2(_3668_),
    .B1(_0067_),
    .C1(_0068_),
    .X(_0069_));
 sky130_fd_sc_hd__a211oi_1 _4697_ (.A1(_0067_),
    .A2(_0068_),
    .B1(_0017_),
    .C1(_3668_),
    .Y(_0070_));
 sky130_fd_sc_hd__or3_2 _4698_ (.A(_0016_),
    .B(_0069_),
    .C(_0070_),
    .X(_0071_));
 sky130_fd_sc_hd__o21ai_2 _4699_ (.A1(_0069_),
    .A2(_0070_),
    .B1(_0016_),
    .Y(_0072_));
 sky130_fd_sc_hd__o211ai_4 _4700_ (.A1(_3670_),
    .A2(_3672_),
    .B1(_0071_),
    .C1(_0072_),
    .Y(_0073_));
 sky130_fd_sc_hd__a211o_1 _4701_ (.A1(_0071_),
    .A2(_0072_),
    .B1(_3670_),
    .C1(_3672_),
    .X(_0075_));
 sky130_fd_sc_hd__nand2_1 _4702_ (.A(_0073_),
    .B(_0075_),
    .Y(_0076_));
 sky130_fd_sc_hd__a21boi_1 _4703_ (.A1(_3612_),
    .A2(_3675_),
    .B1_N(net151),
    .Y(_0077_));
 sky130_fd_sc_hd__xnor2_1 _4704_ (.A(_0076_),
    .B(_0077_),
    .Y(_0078_));
 sky130_fd_sc_hd__nor2_1 _4705_ (.A(_3679_),
    .B(_0078_),
    .Y(_0079_));
 sky130_fd_sc_hd__and2_1 _4706_ (.A(_3679_),
    .B(_0078_),
    .X(_0080_));
 sky130_fd_sc_hd__nor2_1 _4707_ (.A(_0079_),
    .B(_0080_),
    .Y(_0081_));
 sky130_fd_sc_hd__nor2_1 _4708_ (.A(_3610_),
    .B(_3681_),
    .Y(_0082_));
 sky130_fd_sc_hd__a21o_1 _4709_ (.A1(_3609_),
    .A2(_3682_),
    .B1(_0082_),
    .X(_0083_));
 sky130_fd_sc_hd__nor2_1 _4710_ (.A(_0081_),
    .B(net142),
    .Y(_0084_));
 sky130_fd_sc_hd__and2_1 _4711_ (.A(_0081_),
    .B(_0083_),
    .X(_0086_));
 sky130_fd_sc_hd__nor2_1 _4712_ (.A(_0084_),
    .B(_0086_),
    .Y(_0087_));
 sky130_fd_sc_hd__a32o_1 _4713_ (.A1(_0652_),
    .A2(_0013_),
    .A3(_0014_),
    .B1(_0087_),
    .B2(_3305_),
    .X(_0088_));
 sky130_fd_sc_hd__or4_1 _4714_ (.A(_3726_),
    .B(_3732_),
    .C(_0010_),
    .D(_0088_),
    .X(_0089_));
 sky130_fd_sc_hd__buf_6 _4715_ (.A(_0089_),
    .X(net72));
 sky130_fd_sc_hd__nand3_1 _4716_ (.A(_3612_),
    .B(net149),
    .C(_3675_),
    .Y(_0090_));
 sky130_fd_sc_hd__and2b_1 _4717_ (.A_N(_0018_),
    .B(_0027_),
    .X(_0091_));
 sky130_fd_sc_hd__a21oi_2 _4718_ (.A1(_3624_),
    .A2(_0028_),
    .B1(_0091_),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _4719_ (.A(_0065_),
    .Y(_0093_));
 sky130_fd_sc_hd__nand2_1 _4720_ (.A(_0024_),
    .B(_0025_),
    .Y(_0094_));
 sky130_fd_sc_hd__or2b_1 _4721_ (.A(_0019_),
    .B_N(_0026_),
    .X(_0096_));
 sky130_fd_sc_hd__or2b_1 _4722_ (.A(_0033_),
    .B_N(_0038_),
    .X(_0097_));
 sky130_fd_sc_hd__nand2_1 _4723_ (.A(_0032_),
    .B(_0039_),
    .Y(_0098_));
 sky130_fd_sc_hd__clkbuf_4 _4724_ (.A(net37),
    .X(_0099_));
 sky130_fd_sc_hd__clkbuf_4 _4725_ (.A(_0099_),
    .X(_0100_));
 sky130_fd_sc_hd__a22oi_1 _4726_ (.A1(_0707_),
    .A2(_3719_),
    .B1(_0100_),
    .B2(_0477_),
    .Y(_0101_));
 sky130_fd_sc_hd__and4_1 _4727_ (.A(_0707_),
    .B(_0466_),
    .C(_3719_),
    .D(_0100_),
    .X(_0102_));
 sky130_fd_sc_hd__nor2_1 _4728_ (.A(_0101_),
    .B(_0102_),
    .Y(_0103_));
 sky130_fd_sc_hd__clkbuf_4 _4729_ (.A(net64),
    .X(_0104_));
 sky130_fd_sc_hd__clkbuf_4 _4730_ (.A(_3572_),
    .X(_0105_));
 sky130_fd_sc_hd__a22oi_1 _4731_ (.A1(_3440_),
    .A2(_0104_),
    .B1(_0105_),
    .B2(_0194_),
    .Y(_0107_));
 sky130_fd_sc_hd__and4_1 _4732_ (.A(_0085_),
    .B(_0194_),
    .C(_3422_),
    .D(_3511_),
    .X(_0108_));
 sky130_fd_sc_hd__and4bb_1 _4733_ (.A_N(_0107_),
    .B_N(_0108_),
    .C(_0739_),
    .D(_3619_),
    .X(_0109_));
 sky130_fd_sc_hd__clkbuf_4 _4734_ (.A(net35),
    .X(_0110_));
 sky130_fd_sc_hd__o2bb2a_1 _4735_ (.A1_N(_0335_),
    .A2_N(_0110_),
    .B1(_0107_),
    .B2(_0108_),
    .X(_0111_));
 sky130_fd_sc_hd__nor2_1 _4736_ (.A(_0109_),
    .B(_0111_),
    .Y(_0112_));
 sky130_fd_sc_hd__nor2_1 _4737_ (.A(_0021_),
    .B(_0022_),
    .Y(_0113_));
 sky130_fd_sc_hd__xnor2_2 _4738_ (.A(_0112_),
    .B(_0113_),
    .Y(_0114_));
 sky130_fd_sc_hd__xnor2_2 _4739_ (.A(_0103_),
    .B(_0114_),
    .Y(_0115_));
 sky130_fd_sc_hd__a21oi_2 _4740_ (.A1(_0097_),
    .A2(_0098_),
    .B1(_0115_),
    .Y(_0116_));
 sky130_fd_sc_hd__and3_1 _4741_ (.A(_0097_),
    .B(_0098_),
    .C(_0115_),
    .X(_0118_));
 sky130_fd_sc_hd__a211oi_2 _4742_ (.A1(_0094_),
    .A2(_0096_),
    .B1(_0116_),
    .C1(_0118_),
    .Y(_0119_));
 sky130_fd_sc_hd__o211a_1 _4743_ (.A1(_0116_),
    .A2(_0118_),
    .B1(_0094_),
    .C1(_0096_),
    .X(_0120_));
 sky130_fd_sc_hd__nand3_2 _4744_ (.A(_0040_),
    .B(_0060_),
    .C(_0061_),
    .Y(_0121_));
 sky130_fd_sc_hd__a32o_1 _4745_ (.A1(_0106_),
    .A2(_3386_),
    .A3(_0036_),
    .B1(_0035_),
    .B2(_2324_),
    .X(_0122_));
 sky130_fd_sc_hd__o21ba_1 _4746_ (.A1(_0043_),
    .A2(_0044_),
    .B1_N(_0045_),
    .X(_0123_));
 sky130_fd_sc_hd__nand2_1 _4747_ (.A(_2313_),
    .B(_3631_),
    .Y(_0124_));
 sky130_fd_sc_hd__a22o_1 _4748_ (.A1(_3195_),
    .A2(_2423_),
    .B1(_3633_),
    .B2(_2368_),
    .X(_0125_));
 sky130_fd_sc_hd__a21bo_1 _4749_ (.A1(_3530_),
    .A2(_0035_),
    .B1_N(_0125_),
    .X(_0126_));
 sky130_fd_sc_hd__xor2_2 _4750_ (.A(_0124_),
    .B(_0126_),
    .X(_0127_));
 sky130_fd_sc_hd__xnor2_1 _4751_ (.A(_0123_),
    .B(_0127_),
    .Y(_0129_));
 sky130_fd_sc_hd__xor2_1 _4752_ (.A(_0122_),
    .B(_0129_),
    .X(_0130_));
 sky130_fd_sc_hd__nand2_1 _4753_ (.A(_2881_),
    .B(_3644_),
    .Y(_0131_));
 sky130_fd_sc_hd__a22oi_1 _4754_ (.A1(_0041_),
    .A2(_2149_),
    .B1(_2204_),
    .B2(_3645_),
    .Y(_0132_));
 sky130_fd_sc_hd__and4_1 _4755_ (.A(_0161_),
    .B(_3531_),
    .C(net32),
    .D(_3537_),
    .X(_0133_));
 sky130_fd_sc_hd__nor2_1 _4756_ (.A(_0132_),
    .B(_0133_),
    .Y(_0134_));
 sky130_fd_sc_hd__xnor2_2 _4757_ (.A(_0131_),
    .B(_0134_),
    .Y(_0135_));
 sky130_fd_sc_hd__and2_1 _4758_ (.A(_0281_),
    .B(_3651_),
    .X(_0136_));
 sky130_fd_sc_hd__a22o_1 _4759_ (.A1(net178),
    .A2(_2642_),
    .B1(_2686_),
    .B2(_3242_),
    .X(_0137_));
 sky130_fd_sc_hd__nand4_1 _4760_ (.A(_3449_),
    .B(_3448_),
    .C(_2642_),
    .D(_2686_),
    .Y(_0138_));
 sky130_fd_sc_hd__nand3_1 _4761_ (.A(_0136_),
    .B(_0137_),
    .C(_0138_),
    .Y(_0140_));
 sky130_fd_sc_hd__a21o_1 _4762_ (.A1(_0137_),
    .A2(_0138_),
    .B1(_0136_),
    .X(_0141_));
 sky130_fd_sc_hd__a21bo_1 _4763_ (.A1(_0048_),
    .A2(_0049_),
    .B1_N(_0050_),
    .X(_0142_));
 sky130_fd_sc_hd__nand3_1 _4764_ (.A(_0140_),
    .B(_0141_),
    .C(_0142_),
    .Y(_0143_));
 sky130_fd_sc_hd__a21o_1 _4765_ (.A1(_0140_),
    .A2(_0141_),
    .B1(_0142_),
    .X(_0144_));
 sky130_fd_sc_hd__nand3_1 _4766_ (.A(_0135_),
    .B(_0143_),
    .C(_0144_),
    .Y(_0145_));
 sky130_fd_sc_hd__a21o_1 _4767_ (.A1(_0143_),
    .A2(_0144_),
    .B1(_0135_),
    .X(_0146_));
 sky130_fd_sc_hd__a21bo_1 _4768_ (.A1(_0047_),
    .A2(_0056_),
    .B1_N(_0055_),
    .X(_0147_));
 sky130_fd_sc_hd__nand3_2 _4769_ (.A(_0145_),
    .B(_0146_),
    .C(_0147_),
    .Y(_0148_));
 sky130_fd_sc_hd__a21o_1 _4770_ (.A1(_0145_),
    .A2(_0146_),
    .B1(_0147_),
    .X(_0149_));
 sky130_fd_sc_hd__and3_1 _4771_ (.A(_0130_),
    .B(_0148_),
    .C(_0149_),
    .X(_0151_));
 sky130_fd_sc_hd__a21oi_2 _4772_ (.A1(_0148_),
    .A2(_0149_),
    .B1(_0130_),
    .Y(_0152_));
 sky130_fd_sc_hd__a211oi_4 _4773_ (.A1(_0060_),
    .A2(_0121_),
    .B1(_0151_),
    .C1(_0152_),
    .Y(_0153_));
 sky130_fd_sc_hd__o211a_1 _4774_ (.A1(_0151_),
    .A2(_0152_),
    .B1(_0060_),
    .C1(_0121_),
    .X(_0154_));
 sky130_fd_sc_hd__nor4_1 _4775_ (.A(_0119_),
    .B(_0120_),
    .C(_0153_),
    .D(_0154_),
    .Y(_0155_));
 sky130_fd_sc_hd__o22a_1 _4776_ (.A1(_0119_),
    .A2(_0120_),
    .B1(_0153_),
    .B2(_0154_),
    .X(_0156_));
 sky130_fd_sc_hd__a211oi_1 _4777_ (.A1(_0093_),
    .A2(_0067_),
    .B1(net116),
    .C1(_0156_),
    .Y(_0157_));
 sky130_fd_sc_hd__o211a_1 _4778_ (.A1(net116),
    .A2(_0156_),
    .B1(_0093_),
    .C1(_0067_),
    .X(_0158_));
 sky130_fd_sc_hd__nor2_1 _4779_ (.A(_0157_),
    .B(_0158_),
    .Y(_0159_));
 sky130_fd_sc_hd__xnor2_2 _4780_ (.A(_0092_),
    .B(_0159_),
    .Y(_0160_));
 sky130_fd_sc_hd__or2b_1 _4781_ (.A(_0069_),
    .B_N(_0071_),
    .X(_0162_));
 sky130_fd_sc_hd__xnor2_2 _4782_ (.A(_0160_),
    .B(_0162_),
    .Y(_0163_));
 sky130_fd_sc_hd__a211oi_1 _4783_ (.A1(_0071_),
    .A2(_0072_),
    .B1(_3670_),
    .C1(_3672_),
    .Y(_0164_));
 sky130_fd_sc_hd__o21a_1 _4784_ (.A1(_3674_),
    .A2(_0164_),
    .B1(_0073_),
    .X(_0165_));
 sky130_fd_sc_hd__xnor2_1 _4785_ (.A(_0163_),
    .B(_0165_),
    .Y(_0166_));
 sky130_fd_sc_hd__or3_1 _4786_ (.A(_0090_),
    .B(_0076_),
    .C(_0166_),
    .X(_0167_));
 sky130_fd_sc_hd__inv_2 _4787_ (.A(_0167_),
    .Y(_0168_));
 sky130_fd_sc_hd__o21a_1 _4788_ (.A1(_0090_),
    .A2(_0076_),
    .B1(_0166_),
    .X(_0169_));
 sky130_fd_sc_hd__nor2_1 _4789_ (.A(_0168_),
    .B(_0169_),
    .Y(_0170_));
 sky130_fd_sc_hd__o21ai_1 _4790_ (.A1(_0079_),
    .A2(_0086_),
    .B1(_0170_),
    .Y(_0171_));
 sky130_fd_sc_hd__or3_1 _4791_ (.A(_0079_),
    .B(_0086_),
    .C(_0170_),
    .X(_0173_));
 sky130_fd_sc_hd__clkbuf_4 _4792_ (.A(_0100_),
    .X(_0174_));
 sky130_fd_sc_hd__nand2_1 _4793_ (.A(_3133_),
    .B(_0174_),
    .Y(_0175_));
 sky130_fd_sc_hd__or2_1 _4794_ (.A(_2718_),
    .B(_0174_),
    .X(_0176_));
 sky130_fd_sc_hd__nand2_1 _4795_ (.A(_0175_),
    .B(_0176_),
    .Y(_0177_));
 sky130_fd_sc_hd__inv_2 _4796_ (.A(_2664_),
    .Y(_0178_));
 sky130_fd_sc_hd__nor2_1 _4797_ (.A(_0178_),
    .B(_3720_),
    .Y(_0179_));
 sky130_fd_sc_hd__a21o_1 _4798_ (.A1(_3723_),
    .A2(_0012_),
    .B1(_0179_),
    .X(_0180_));
 sky130_fd_sc_hd__clkbuf_4 _4799_ (.A(_3265_),
    .X(_0181_));
 sky130_fd_sc_hd__a21oi_1 _4800_ (.A1(_0177_),
    .A2(_0180_),
    .B1(_0181_),
    .Y(_0182_));
 sky130_fd_sc_hd__o21a_1 _4801_ (.A1(_0177_),
    .A2(_0180_),
    .B1(_0182_),
    .X(_0184_));
 sky130_fd_sc_hd__or3b_1 _4802_ (.A(_3722_),
    .B(_3724_),
    .C_N(_0177_),
    .X(_0185_));
 sky130_fd_sc_hd__o21bai_1 _4803_ (.A1(_3722_),
    .A2(_3724_),
    .B1_N(_0177_),
    .Y(_0186_));
 sky130_fd_sc_hd__mux4_2 _4804_ (.A0(_3133_),
    .A1(_2675_),
    .A2(_3137_),
    .A3(_2237_),
    .S0(_3046_),
    .S1(_3591_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _4805_ (.A0(_3500_),
    .A1(_0187_),
    .S(_3087_),
    .X(_0188_));
 sky130_fd_sc_hd__clkbuf_4 _4806_ (.A(_3301_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _4807_ (.A0(_3097_),
    .A1(_0188_),
    .S(_0189_),
    .X(_0190_));
 sky130_fd_sc_hd__and2_1 _4808_ (.A(_2707_),
    .B(_0100_),
    .X(_0191_));
 sky130_fd_sc_hd__inv_2 _4809_ (.A(_0176_),
    .Y(_0192_));
 sky130_fd_sc_hd__a21o_1 _4810_ (.A1(net124),
    .A2(_0175_),
    .B1(_3204_),
    .X(_0193_));
 sky130_fd_sc_hd__or3_1 _4811_ (.A(_0980_),
    .B(_0870_),
    .C(_0969_),
    .X(_0195_));
 sky130_fd_sc_hd__buf_2 _4812_ (.A(_0195_),
    .X(_0196_));
 sky130_fd_sc_hd__a22o_1 _4813_ (.A1(_0176_),
    .A2(_0193_),
    .B1(_0196_),
    .B2(_3201_),
    .X(_0197_));
 sky130_fd_sc_hd__a221o_1 _4814_ (.A1(_3194_),
    .A2(_0191_),
    .B1(_0192_),
    .B2(_3414_),
    .C1(_0197_),
    .X(_0198_));
 sky130_fd_sc_hd__clkbuf_4 _4815_ (.A(_3486_),
    .X(_0199_));
 sky130_fd_sc_hd__mux4_1 _4816_ (.A0(_3132_),
    .A1(_3136_),
    .A2(_3148_),
    .A3(_3151_),
    .S0(_3087_),
    .S1(_0199_),
    .X(_0200_));
 sky130_fd_sc_hd__or3_1 _4817_ (.A(_3490_),
    .B(_3486_),
    .C(_3145_),
    .X(_0201_));
 sky130_fd_sc_hd__nand2_1 _4818_ (.A(_3580_),
    .B(_0201_),
    .Y(_0202_));
 sky130_fd_sc_hd__o211a_1 _4819_ (.A1(_3580_),
    .A2(_0200_),
    .B1(_0202_),
    .C1(_3587_),
    .X(_0203_));
 sky130_fd_sc_hd__a211o_1 _4820_ (.A1(_0007_),
    .A2(_0190_),
    .B1(_0198_),
    .C1(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__a31o_1 _4821_ (.A1(_2980_),
    .A2(_0185_),
    .A3(_0186_),
    .B1(_0204_),
    .X(_0206_));
 sky130_fd_sc_hd__a311o_4 _4822_ (.A1(_3305_),
    .A2(_0171_),
    .A3(_0173_),
    .B1(_0184_),
    .C1(_0206_),
    .X(net73));
 sky130_fd_sc_hd__or3_1 _4823_ (.A(net150),
    .B(_0076_),
    .C(_0163_),
    .X(_0207_));
 sky130_fd_sc_hd__o21ai_1 _4824_ (.A1(_0116_),
    .A2(_0119_),
    .B1(_0102_),
    .Y(_0208_));
 sky130_fd_sc_hd__or3_1 _4825_ (.A(_0102_),
    .B(_0116_),
    .C(_0119_),
    .X(_0209_));
 sky130_fd_sc_hd__and2_1 _4826_ (.A(_0208_),
    .B(_0209_),
    .X(_0210_));
 sky130_fd_sc_hd__nand2_1 _4827_ (.A(_0103_),
    .B(_0114_),
    .Y(_0211_));
 sky130_fd_sc_hd__o31a_1 _4828_ (.A1(_0109_),
    .A2(_0111_),
    .A3(_0113_),
    .B1(_0211_),
    .X(_0212_));
 sky130_fd_sc_hd__and2b_1 _4829_ (.A_N(_0123_),
    .B(_0127_),
    .X(_0213_));
 sky130_fd_sc_hd__and2_1 _4830_ (.A(_0122_),
    .B(_0129_),
    .X(_0214_));
 sky130_fd_sc_hd__a22oi_1 _4831_ (.A1(_0335_),
    .A2(_3718_),
    .B1(_0100_),
    .B2(_0423_),
    .Y(_0216_));
 sky130_fd_sc_hd__and4_1 _4832_ (.A(_0739_),
    .B(_0423_),
    .C(_3718_),
    .D(_0099_),
    .X(_0217_));
 sky130_fd_sc_hd__nor2_1 _4833_ (.A(_0216_),
    .B(_0217_),
    .Y(_0218_));
 sky130_fd_sc_hd__clkbuf_4 _4834_ (.A(net38),
    .X(_0219_));
 sky130_fd_sc_hd__clkbuf_4 _4835_ (.A(_0219_),
    .X(_0220_));
 sky130_fd_sc_hd__nand2_1 _4836_ (.A(_0466_),
    .B(_0220_),
    .Y(_0221_));
 sky130_fd_sc_hd__xor2_2 _4837_ (.A(_0218_),
    .B(_0221_),
    .X(_0222_));
 sky130_fd_sc_hd__a22oi_1 _4838_ (.A1(_3635_),
    .A2(_0104_),
    .B1(_0105_),
    .B2(_3440_),
    .Y(_0223_));
 sky130_fd_sc_hd__and4_1 _4839_ (.A(_0085_),
    .B(_2302_),
    .C(_3422_),
    .D(_3572_),
    .X(_0224_));
 sky130_fd_sc_hd__and4bb_1 _4840_ (.A_N(_0223_),
    .B_N(_0224_),
    .C(_1275_),
    .D(_3619_),
    .X(_0225_));
 sky130_fd_sc_hd__o2bb2a_1 _4841_ (.A1_N(_0205_),
    .A2_N(_0110_),
    .B1(_0223_),
    .B2(_0224_),
    .X(_0227_));
 sky130_fd_sc_hd__nor2_1 _4842_ (.A(_0225_),
    .B(_0227_),
    .Y(_0228_));
 sky130_fd_sc_hd__nor2_1 _4843_ (.A(_0108_),
    .B(_0109_),
    .Y(_0229_));
 sky130_fd_sc_hd__xnor2_1 _4844_ (.A(_0228_),
    .B(_0229_),
    .Y(_0230_));
 sky130_fd_sc_hd__xnor2_1 _4845_ (.A(_0222_),
    .B(_0230_),
    .Y(_0231_));
 sky130_fd_sc_hd__o21a_1 _4846_ (.A1(_0213_),
    .A2(_0214_),
    .B1(_0231_),
    .X(_0232_));
 sky130_fd_sc_hd__nor3_1 _4847_ (.A(_0213_),
    .B(_0214_),
    .C(_0231_),
    .Y(_0233_));
 sky130_fd_sc_hd__nor3_1 _4848_ (.A(_0212_),
    .B(_0232_),
    .C(_0233_),
    .Y(_0234_));
 sky130_fd_sc_hd__o21a_1 _4849_ (.A1(_0232_),
    .A2(_0233_),
    .B1(_0212_),
    .X(_0235_));
 sky130_fd_sc_hd__nand3_1 _4850_ (.A(_0130_),
    .B(_0148_),
    .C(_0149_),
    .Y(_0236_));
 sky130_fd_sc_hd__a32o_1 _4851_ (.A1(_2324_),
    .A2(_3385_),
    .A3(_0125_),
    .B1(_0035_),
    .B2(_2445_),
    .X(_0238_));
 sky130_fd_sc_hd__o21ba_1 _4852_ (.A1(_0131_),
    .A2(_0132_),
    .B1_N(_0133_),
    .X(_0239_));
 sky130_fd_sc_hd__nand2_1 _4853_ (.A(_2379_),
    .B(_3430_),
    .Y(_0240_));
 sky130_fd_sc_hd__and3_1 _4854_ (.A(_2423_),
    .B(net162),
    .C(net31),
    .X(_0241_));
 sky130_fd_sc_hd__a22o_1 _4855_ (.A1(_2423_),
    .A2(net162),
    .B1(net31),
    .B2(_3433_),
    .X(_0242_));
 sky130_fd_sc_hd__a21bo_1 _4856_ (.A1(_3632_),
    .A2(_0241_),
    .B1_N(_0242_),
    .X(_0243_));
 sky130_fd_sc_hd__xor2_2 _4857_ (.A(_0240_),
    .B(_0243_),
    .X(_0244_));
 sky130_fd_sc_hd__xnor2_1 _4858_ (.A(_0239_),
    .B(_0244_),
    .Y(_0245_));
 sky130_fd_sc_hd__xor2_1 _4859_ (.A(_0238_),
    .B(_0245_),
    .X(_0246_));
 sky130_fd_sc_hd__clkbuf_4 _4860_ (.A(net32),
    .X(_0247_));
 sky130_fd_sc_hd__nand2_1 _4861_ (.A(_2881_),
    .B(_0247_),
    .Y(_0249_));
 sky130_fd_sc_hd__a22oi_2 _4862_ (.A1(_3531_),
    .A2(_3537_),
    .B1(_2248_),
    .B2(_3645_),
    .Y(_0250_));
 sky130_fd_sc_hd__and4_1 _4863_ (.A(_0161_),
    .B(_3531_),
    .C(_3537_),
    .D(_3651_),
    .X(_0251_));
 sky130_fd_sc_hd__nor2_1 _4864_ (.A(_0250_),
    .B(_0251_),
    .Y(_0252_));
 sky130_fd_sc_hd__xnor2_2 _4865_ (.A(_0249_),
    .B(_0252_),
    .Y(_0253_));
 sky130_fd_sc_hd__and2_1 _4866_ (.A(_0281_),
    .B(_2642_),
    .X(_0254_));
 sky130_fd_sc_hd__a22o_1 _4867_ (.A1(net178),
    .A2(net5),
    .B1(net6),
    .B2(_3242_),
    .X(_0255_));
 sky130_fd_sc_hd__nand4_1 _4868_ (.A(_3449_),
    .B(_3448_),
    .C(_2686_),
    .D(net6),
    .Y(_0256_));
 sky130_fd_sc_hd__nand3_1 _4869_ (.A(_0254_),
    .B(_0255_),
    .C(_0256_),
    .Y(_0257_));
 sky130_fd_sc_hd__a21o_1 _4870_ (.A1(_0255_),
    .A2(_0256_),
    .B1(_0254_),
    .X(_0258_));
 sky130_fd_sc_hd__a21bo_1 _4871_ (.A1(_0136_),
    .A2(_0137_),
    .B1_N(_0138_),
    .X(_0260_));
 sky130_fd_sc_hd__nand3_1 _4872_ (.A(_0257_),
    .B(_0258_),
    .C(_0260_),
    .Y(_0261_));
 sky130_fd_sc_hd__a21o_1 _4873_ (.A1(_0257_),
    .A2(_0258_),
    .B1(_0260_),
    .X(_0262_));
 sky130_fd_sc_hd__nand3_1 _4874_ (.A(_0253_),
    .B(_0261_),
    .C(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__a21o_1 _4875_ (.A1(_0261_),
    .A2(_0262_),
    .B1(_0253_),
    .X(_0264_));
 sky130_fd_sc_hd__a21bo_1 _4876_ (.A1(_0135_),
    .A2(_0144_),
    .B1_N(_0143_),
    .X(_0265_));
 sky130_fd_sc_hd__nand3_2 _4877_ (.A(_0263_),
    .B(_0264_),
    .C(_0265_),
    .Y(_0266_));
 sky130_fd_sc_hd__a21o_1 _4878_ (.A1(_0263_),
    .A2(_0264_),
    .B1(_0265_),
    .X(_0267_));
 sky130_fd_sc_hd__and3_1 _4879_ (.A(_0246_),
    .B(_0266_),
    .C(_0267_),
    .X(_0268_));
 sky130_fd_sc_hd__a21oi_1 _4880_ (.A1(_0266_),
    .A2(_0267_),
    .B1(_0246_),
    .Y(_0269_));
 sky130_fd_sc_hd__a211o_1 _4881_ (.A1(_0148_),
    .A2(_0236_),
    .B1(_0268_),
    .C1(_0269_),
    .X(_0271_));
 sky130_fd_sc_hd__o211ai_1 _4882_ (.A1(_0268_),
    .A2(_0269_),
    .B1(_0148_),
    .C1(_0236_),
    .Y(_0272_));
 sky130_fd_sc_hd__or4bb_4 _4883_ (.A(_0234_),
    .B(_0235_),
    .C_N(_0271_),
    .D_N(_0272_),
    .X(_0273_));
 sky130_fd_sc_hd__a2bb2o_1 _4884_ (.A1_N(_0234_),
    .A2_N(_0235_),
    .B1(_0271_),
    .B2(_0272_),
    .X(_0274_));
 sky130_fd_sc_hd__o211ai_2 _4885_ (.A1(_0153_),
    .A2(net116),
    .B1(_0273_),
    .C1(_0274_),
    .Y(_0275_));
 sky130_fd_sc_hd__a211o_1 _4886_ (.A1(_0273_),
    .A2(_0274_),
    .B1(_0153_),
    .C1(_0155_),
    .X(_0276_));
 sky130_fd_sc_hd__and3_1 _4887_ (.A(_0210_),
    .B(_0275_),
    .C(_0276_),
    .X(_0277_));
 sky130_fd_sc_hd__a21oi_1 _4888_ (.A1(_0275_),
    .A2(_0276_),
    .B1(_0210_),
    .Y(_0278_));
 sky130_fd_sc_hd__nor2_2 _4889_ (.A(_0277_),
    .B(_0278_),
    .Y(_0279_));
 sky130_fd_sc_hd__o21bai_2 _4890_ (.A1(_0092_),
    .A2(_0158_),
    .B1_N(_0157_),
    .Y(_0280_));
 sky130_fd_sc_hd__xnor2_2 _4891_ (.A(_0279_),
    .B(_0280_),
    .Y(_0282_));
 sky130_fd_sc_hd__nand2_1 _4892_ (.A(_0160_),
    .B(_0162_),
    .Y(_0283_));
 sky130_fd_sc_hd__o21a_1 _4893_ (.A1(_0073_),
    .A2(_0163_),
    .B1(_0283_),
    .X(_0284_));
 sky130_fd_sc_hd__xnor2_1 _4894_ (.A(_0282_),
    .B(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__xnor2_1 _4895_ (.A(_0207_),
    .B(_0285_),
    .Y(_0286_));
 sky130_fd_sc_hd__inv_2 _4896_ (.A(_0286_),
    .Y(_0287_));
 sky130_fd_sc_hd__o21bai_1 _4897_ (.A1(_0079_),
    .A2(_0168_),
    .B1_N(_0169_),
    .Y(_0288_));
 sky130_fd_sc_hd__a21bo_1 _4898_ (.A1(_0086_),
    .A2(_0170_),
    .B1_N(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__nor2_1 _4899_ (.A(_0287_),
    .B(_0289_),
    .Y(_0290_));
 sky130_fd_sc_hd__a21o_1 _4900_ (.A1(_0287_),
    .A2(_0289_),
    .B1(_3192_),
    .X(_0291_));
 sky130_fd_sc_hd__clkbuf_4 _4901_ (.A(_0220_),
    .X(_0293_));
 sky130_fd_sc_hd__or2_1 _4902_ (.A(_3134_),
    .B(_0293_),
    .X(_0294_));
 sky130_fd_sc_hd__nand2_2 _4903_ (.A(_2762_),
    .B(_0293_),
    .Y(_0295_));
 sky130_fd_sc_hd__nand2_1 _4904_ (.A(_0294_),
    .B(_0295_),
    .Y(_0296_));
 sky130_fd_sc_hd__and2b_1 _4905_ (.A_N(_0174_),
    .B(_3133_),
    .X(_0297_));
 sky130_fd_sc_hd__a21o_1 _4906_ (.A1(_0177_),
    .A2(_0180_),
    .B1(_0297_),
    .X(_0298_));
 sky130_fd_sc_hd__nor2_1 _4907_ (.A(_0296_),
    .B(_0298_),
    .Y(_0299_));
 sky130_fd_sc_hd__and2_1 _4908_ (.A(_0296_),
    .B(_0298_),
    .X(_0300_));
 sky130_fd_sc_hd__a21o_1 _4909_ (.A1(_0175_),
    .A2(_0186_),
    .B1(_0296_),
    .X(_0301_));
 sky130_fd_sc_hd__a31oi_1 _4910_ (.A1(_0175_),
    .A2(_0186_),
    .A3(_0296_),
    .B1(_3596_),
    .Y(_0302_));
 sky130_fd_sc_hd__mux4_2 _4911_ (.A0(_3134_),
    .A1(_3133_),
    .A2(_2675_),
    .A3(_3137_),
    .S0(_3046_),
    .S1(_3591_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _4912_ (.A0(_3602_),
    .A1(_0304_),
    .S(_3087_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _4913_ (.A0(_3213_),
    .A1(_0305_),
    .S(_3301_),
    .X(_0306_));
 sky130_fd_sc_hd__a21o_1 _4914_ (.A1(net124),
    .A2(_0295_),
    .B1(_3204_),
    .X(_0307_));
 sky130_fd_sc_hd__or4b_1 _4915_ (.A(net65),
    .B(_1144_),
    .C(_1154_),
    .D_N(_1165_),
    .X(_0308_));
 sky130_fd_sc_hd__clkbuf_4 _4916_ (.A(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__o22ai_1 _4917_ (.A1(_3712_),
    .A2(_0294_),
    .B1(_0295_),
    .B2(_0309_),
    .Y(_0310_));
 sky130_fd_sc_hd__a221o_1 _4918_ (.A1(_3201_),
    .A2(_0196_),
    .B1(_0294_),
    .B2(_0307_),
    .C1(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__mux4_1 _4919_ (.A0(_3219_),
    .A1(_3220_),
    .A2(_3224_),
    .A3(_3225_),
    .S0(_3087_),
    .S1(_3486_),
    .X(_0312_));
 sky130_fd_sc_hd__or2b_1 _4920_ (.A(_0196_),
    .B_N(_2062_),
    .X(_0313_));
 sky130_fd_sc_hd__nand2_1 _4921_ (.A(_3580_),
    .B(_0313_),
    .Y(_0315_));
 sky130_fd_sc_hd__o211a_1 _4922_ (.A1(_3580_),
    .A2(_0312_),
    .B1(_0315_),
    .C1(_3587_),
    .X(_0316_));
 sky130_fd_sc_hd__a211o_1 _4923_ (.A1(_0007_),
    .A2(_0306_),
    .B1(_0311_),
    .C1(_0316_),
    .X(_0317_));
 sky130_fd_sc_hd__a21oi_1 _4924_ (.A1(_0301_),
    .A2(_0302_),
    .B1(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hd__o31a_2 _4925_ (.A1(_0181_),
    .A2(_0299_),
    .A3(_0300_),
    .B1(_0318_),
    .X(_0319_));
 sky130_fd_sc_hd__o21ai_4 _4926_ (.A1(_0290_),
    .A2(_0291_),
    .B1(_0319_),
    .Y(net74));
 sky130_fd_sc_hd__clkbuf_4 _4927_ (.A(_3305_),
    .X(_0320_));
 sky130_fd_sc_hd__nor3_1 _4928_ (.A(_0073_),
    .B(_0163_),
    .C(_0282_),
    .Y(_0321_));
 sky130_fd_sc_hd__or2_2 _4929_ (.A(_0232_),
    .B(_0234_),
    .X(_0322_));
 sky130_fd_sc_hd__a31o_1 _4930_ (.A1(_1002_),
    .A2(_0293_),
    .A3(_0218_),
    .B1(_0217_),
    .X(_0323_));
 sky130_fd_sc_hd__buf_2 _4931_ (.A(net39),
    .X(_0325_));
 sky130_fd_sc_hd__buf_2 _4932_ (.A(_0325_),
    .X(_0326_));
 sky130_fd_sc_hd__buf_2 _4933_ (.A(_0326_),
    .X(_0327_));
 sky130_fd_sc_hd__clkbuf_4 _4934_ (.A(_0327_),
    .X(_0328_));
 sky130_fd_sc_hd__nand2_1 _4935_ (.A(_1384_),
    .B(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__xnor2_2 _4936_ (.A(_0323_),
    .B(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__xnor2_2 _4937_ (.A(_0322_),
    .B(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hd__or3_2 _4938_ (.A(_0225_),
    .B(_0227_),
    .C(_0229_),
    .X(_0332_));
 sky130_fd_sc_hd__or2b_1 _4939_ (.A(_0222_),
    .B_N(_0230_),
    .X(_0333_));
 sky130_fd_sc_hd__and2b_1 _4940_ (.A_N(_0239_),
    .B(_0244_),
    .X(_0334_));
 sky130_fd_sc_hd__and2_1 _4941_ (.A(_0238_),
    .B(_0245_),
    .X(_0336_));
 sky130_fd_sc_hd__inv_2 _4942_ (.A(net38),
    .Y(_0337_));
 sky130_fd_sc_hd__a22oi_1 _4943_ (.A1(_0205_),
    .A2(_3718_),
    .B1(_0099_),
    .B2(_0335_),
    .Y(_0338_));
 sky130_fd_sc_hd__clkbuf_8 _4944_ (.A(net36),
    .X(_0339_));
 sky130_fd_sc_hd__buf_4 _4945_ (.A(net37),
    .X(_0340_));
 sky130_fd_sc_hd__and4_1 _4946_ (.A(_1275_),
    .B(_0739_),
    .C(_0339_),
    .D(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__o22a_1 _4947_ (.A1(_1428_),
    .A2(_0337_),
    .B1(_0338_),
    .B2(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__and4bb_1 _4948_ (.A_N(_0338_),
    .B_N(_0341_),
    .C(_0434_),
    .D(_0219_),
    .X(_0343_));
 sky130_fd_sc_hd__or2_1 _4949_ (.A(_0342_),
    .B(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__nand2_1 _4950_ (.A(_0095_),
    .B(_0110_),
    .Y(_0345_));
 sky130_fd_sc_hd__and3_1 _4951_ (.A(_2302_),
    .B(_2368_),
    .C(_3511_),
    .X(_0347_));
 sky130_fd_sc_hd__a22o_1 _4952_ (.A1(_3442_),
    .A2(_3422_),
    .B1(_3511_),
    .B2(_2302_),
    .X(_0348_));
 sky130_fd_sc_hd__a21bo_1 _4953_ (.A1(_3423_),
    .A2(_0347_),
    .B1_N(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__xor2_2 _4954_ (.A(_0345_),
    .B(_0349_),
    .X(_0350_));
 sky130_fd_sc_hd__nor2_1 _4955_ (.A(_0224_),
    .B(_0225_),
    .Y(_0351_));
 sky130_fd_sc_hd__xnor2_1 _4956_ (.A(_0350_),
    .B(_0351_),
    .Y(_0352_));
 sky130_fd_sc_hd__xnor2_1 _4957_ (.A(_0344_),
    .B(_0352_),
    .Y(_0353_));
 sky130_fd_sc_hd__o21a_1 _4958_ (.A1(_0334_),
    .A2(_0336_),
    .B1(_0353_),
    .X(_0354_));
 sky130_fd_sc_hd__nor3_1 _4959_ (.A(_0334_),
    .B(_0336_),
    .C(_0353_),
    .Y(_0355_));
 sky130_fd_sc_hd__a211oi_2 _4960_ (.A1(_0332_),
    .A2(_0333_),
    .B1(_0354_),
    .C1(_0355_),
    .Y(_0356_));
 sky130_fd_sc_hd__o211a_1 _4961_ (.A1(_0354_),
    .A2(_0355_),
    .B1(_0332_),
    .C1(_0333_),
    .X(_0358_));
 sky130_fd_sc_hd__nand3_1 _4962_ (.A(_0246_),
    .B(_0266_),
    .C(net190),
    .Y(_0359_));
 sky130_fd_sc_hd__a32o_1 _4963_ (.A1(_2390_),
    .A2(_3385_),
    .A3(_0242_),
    .B1(_0241_),
    .B2(_3197_),
    .X(_0360_));
 sky130_fd_sc_hd__o21bai_1 _4964_ (.A1(_0249_),
    .A2(_0250_),
    .B1_N(_0251_),
    .Y(_0361_));
 sky130_fd_sc_hd__a22o_1 _4965_ (.A1(_3271_),
    .A2(_2106_),
    .B1(_2149_),
    .B2(_3632_),
    .X(_0362_));
 sky130_fd_sc_hd__nand4_2 _4966_ (.A(_3196_),
    .B(_3271_),
    .C(_3644_),
    .D(_0247_),
    .Y(_0363_));
 sky130_fd_sc_hd__nand4_2 _4967_ (.A(_2445_),
    .B(_3385_),
    .C(_0362_),
    .D(_0363_),
    .Y(_0364_));
 sky130_fd_sc_hd__a22o_1 _4968_ (.A1(_3530_),
    .A2(_3385_),
    .B1(_0362_),
    .B2(_0363_),
    .X(_0365_));
 sky130_fd_sc_hd__nand3_1 _4969_ (.A(_0361_),
    .B(_0364_),
    .C(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__a21o_1 _4970_ (.A1(_0364_),
    .A2(_0365_),
    .B1(_0361_),
    .X(_0367_));
 sky130_fd_sc_hd__and3_1 _4971_ (.A(_0360_),
    .B(_0366_),
    .C(_0367_),
    .X(_0369_));
 sky130_fd_sc_hd__a21oi_1 _4972_ (.A1(_0366_),
    .A2(_0367_),
    .B1(_0360_),
    .Y(_0370_));
 sky130_fd_sc_hd__nor2_1 _4973_ (.A(_0369_),
    .B(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__nand2_1 _4974_ (.A(_0042_),
    .B(_2215_),
    .Y(_0372_));
 sky130_fd_sc_hd__clkbuf_4 _4975_ (.A(net59),
    .X(_0373_));
 sky130_fd_sc_hd__and3_1 _4976_ (.A(_3352_),
    .B(_0373_),
    .C(net3),
    .X(_0374_));
 sky130_fd_sc_hd__a22o_1 _4977_ (.A1(net191),
    .A2(net3),
    .B1(_2642_),
    .B2(_3169_),
    .X(_0375_));
 sky130_fd_sc_hd__a21bo_1 _4978_ (.A1(_2653_),
    .A2(_0374_),
    .B1_N(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__xor2_2 _4979_ (.A(_0372_),
    .B(_0376_),
    .X(_0377_));
 sky130_fd_sc_hd__and2_1 _4980_ (.A(_0292_),
    .B(_2686_),
    .X(_0378_));
 sky130_fd_sc_hd__clkbuf_4 _4981_ (.A(net7),
    .X(_0380_));
 sky130_fd_sc_hd__a22o_1 _4982_ (.A1(_3448_),
    .A2(_2740_),
    .B1(_0380_),
    .B2(_3449_),
    .X(_0381_));
 sky130_fd_sc_hd__nand4_1 _4983_ (.A(_3451_),
    .B(_3452_),
    .C(_2740_),
    .D(_0380_),
    .Y(_0382_));
 sky130_fd_sc_hd__nand3_1 _4984_ (.A(_0378_),
    .B(_0381_),
    .C(_0382_),
    .Y(_0383_));
 sky130_fd_sc_hd__a21o_1 _4985_ (.A1(_0381_),
    .A2(_0382_),
    .B1(_0378_),
    .X(_0384_));
 sky130_fd_sc_hd__a21bo_1 _4986_ (.A1(_0254_),
    .A2(_0255_),
    .B1_N(_0256_),
    .X(_0385_));
 sky130_fd_sc_hd__nand3_1 _4987_ (.A(_0383_),
    .B(_0384_),
    .C(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__a21o_1 _4988_ (.A1(_0383_),
    .A2(_0384_),
    .B1(_0385_),
    .X(_0387_));
 sky130_fd_sc_hd__nand3_1 _4989_ (.A(_0377_),
    .B(_0386_),
    .C(_0387_),
    .Y(_0388_));
 sky130_fd_sc_hd__a21o_1 _4990_ (.A1(_0386_),
    .A2(_0387_),
    .B1(_0377_),
    .X(_0389_));
 sky130_fd_sc_hd__a21bo_1 _4991_ (.A1(_0253_),
    .A2(_0262_),
    .B1_N(_0261_),
    .X(_0391_));
 sky130_fd_sc_hd__nand3_2 _4992_ (.A(_0388_),
    .B(_0389_),
    .C(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__a21o_1 _4993_ (.A1(_0388_),
    .A2(_0389_),
    .B1(_0391_),
    .X(_0393_));
 sky130_fd_sc_hd__and3_1 _4994_ (.A(_0371_),
    .B(_0392_),
    .C(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__a21oi_1 _4995_ (.A1(_0392_),
    .A2(_0393_),
    .B1(_0371_),
    .Y(_0395_));
 sky130_fd_sc_hd__a211oi_2 _4996_ (.A1(_0266_),
    .A2(_0359_),
    .B1(_0394_),
    .C1(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__o211a_1 _4997_ (.A1(_0394_),
    .A2(_0395_),
    .B1(_0266_),
    .C1(_0359_),
    .X(_0397_));
 sky130_fd_sc_hd__nor4_1 _4998_ (.A(_0356_),
    .B(_0358_),
    .C(_0396_),
    .D(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__o22a_1 _4999_ (.A1(_0356_),
    .A2(_0358_),
    .B1(_0396_),
    .B2(_0397_),
    .X(_0399_));
 sky130_fd_sc_hd__a211oi_4 _5000_ (.A1(net156),
    .A2(_0273_),
    .B1(net172),
    .C1(_0399_),
    .Y(_0400_));
 sky130_fd_sc_hd__o211a_1 _5001_ (.A1(net115),
    .A2(_0399_),
    .B1(net156),
    .C1(_0273_),
    .X(_0402_));
 sky130_fd_sc_hd__or3_1 _5002_ (.A(_0331_),
    .B(_0400_),
    .C(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__o21ai_2 _5003_ (.A1(_0400_),
    .A2(_0402_),
    .B1(_0331_),
    .Y(_0404_));
 sky130_fd_sc_hd__a21bo_1 _5004_ (.A1(_0210_),
    .A2(_0276_),
    .B1_N(_0275_),
    .X(_0405_));
 sky130_fd_sc_hd__and3_1 _5005_ (.A(_0403_),
    .B(_0404_),
    .C(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__a21oi_1 _5006_ (.A1(_0403_),
    .A2(_0404_),
    .B1(net179),
    .Y(_0407_));
 sky130_fd_sc_hd__or3_4 _5007_ (.A(_0208_),
    .B(_0406_),
    .C(_0407_),
    .X(_0408_));
 sky130_fd_sc_hd__o21ai_1 _5008_ (.A1(_0406_),
    .A2(_0407_),
    .B1(_0208_),
    .Y(_0409_));
 sky130_fd_sc_hd__nand2_1 _5009_ (.A(net180),
    .B(_0409_),
    .Y(_0410_));
 sky130_fd_sc_hd__nand2_1 _5010_ (.A(_0279_),
    .B(_0280_),
    .Y(_0411_));
 sky130_fd_sc_hd__o21ai_1 _5011_ (.A1(_0283_),
    .A2(_0282_),
    .B1(_0411_),
    .Y(_0413_));
 sky130_fd_sc_hd__xnor2_1 _5012_ (.A(_0410_),
    .B(_0413_),
    .Y(_0414_));
 sky130_fd_sc_hd__xnor2_1 _5013_ (.A(_0321_),
    .B(_0414_),
    .Y(_0415_));
 sky130_fd_sc_hd__nor2_1 _5014_ (.A(_0207_),
    .B(_0285_),
    .Y(_0416_));
 sky130_fd_sc_hd__a21o_1 _5015_ (.A1(_0287_),
    .A2(_0289_),
    .B1(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__xnor2_1 _5016_ (.A(_0415_),
    .B(_0417_),
    .Y(_0418_));
 sky130_fd_sc_hd__clkbuf_4 _5017_ (.A(_2980_),
    .X(_0419_));
 sky130_fd_sc_hd__and2_2 _5018_ (.A(_2784_),
    .B(_0327_),
    .X(_0420_));
 sky130_fd_sc_hd__nor2_1 _5019_ (.A(_3135_),
    .B(_0328_),
    .Y(_0421_));
 sky130_fd_sc_hd__or2_2 _5020_ (.A(_0420_),
    .B(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__nand3_1 _5021_ (.A(_0295_),
    .B(_0301_),
    .C(_0422_),
    .Y(_0424_));
 sky130_fd_sc_hd__a21o_1 _5022_ (.A1(_0295_),
    .A2(_0301_),
    .B1(_0422_),
    .X(_0425_));
 sky130_fd_sc_hd__a21oi_1 _5023_ (.A1(_3134_),
    .A2(_0337_),
    .B1(_0300_),
    .Y(_0426_));
 sky130_fd_sc_hd__xnor2_1 _5024_ (.A(_0422_),
    .B(_0426_),
    .Y(_0427_));
 sky130_fd_sc_hd__buf_2 _5025_ (.A(_3727_),
    .X(_0428_));
 sky130_fd_sc_hd__clkbuf_4 _5026_ (.A(_3087_),
    .X(_0429_));
 sky130_fd_sc_hd__mux4_1 _5027_ (.A0(_3296_),
    .A1(_3298_),
    .A2(_3291_),
    .A3(_3292_),
    .S0(_0429_),
    .S1(_0199_),
    .X(_0430_));
 sky130_fd_sc_hd__o21ai_1 _5028_ (.A1(_3144_),
    .A2(_0196_),
    .B1(_3727_),
    .Y(_0431_));
 sky130_fd_sc_hd__o211a_1 _5029_ (.A1(_0428_),
    .A2(_0430_),
    .B1(_0431_),
    .C1(_3587_),
    .X(_0432_));
 sky130_fd_sc_hd__mux4_2 _5030_ (.A0(_3135_),
    .A1(_3134_),
    .A2(_3133_),
    .A3(_2675_),
    .S0(_3046_),
    .S1(_3591_),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _5031_ (.A0(_3702_),
    .A1(_0433_),
    .S(_0429_),
    .X(_0435_));
 sky130_fd_sc_hd__mux2_1 _5032_ (.A0(_3285_),
    .A1(_0435_),
    .S(_0189_),
    .X(_0436_));
 sky130_fd_sc_hd__a221o_1 _5033_ (.A1(_3194_),
    .A2(_0420_),
    .B1(_0421_),
    .B2(_3414_),
    .C1(_3201_),
    .X(_0437_));
 sky130_fd_sc_hd__clkbuf_4 _5034_ (.A(net124),
    .X(_0438_));
 sky130_fd_sc_hd__nand2_1 _5035_ (.A(_3135_),
    .B(_0328_),
    .Y(_0439_));
 sky130_fd_sc_hd__a21oi_1 _5036_ (.A1(_0438_),
    .A2(_0439_),
    .B1(_0000_),
    .Y(_0440_));
 sky130_fd_sc_hd__nor2_1 _5037_ (.A(_0421_),
    .B(_0440_),
    .Y(_0441_));
 sky130_fd_sc_hd__a211o_1 _5038_ (.A1(_0007_),
    .A2(_0436_),
    .B1(_0437_),
    .C1(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__a211o_1 _5039_ (.A1(_3571_),
    .A2(_0427_),
    .B1(_0432_),
    .C1(_0442_),
    .X(_0443_));
 sky130_fd_sc_hd__a31o_1 _5040_ (.A1(_0419_),
    .A2(_0424_),
    .A3(_0425_),
    .B1(_0443_),
    .X(_0444_));
 sky130_fd_sc_hd__a21o_2 _5041_ (.A1(_0320_),
    .A2(_0418_),
    .B1(_0444_),
    .X(net75));
 sky130_fd_sc_hd__and3b_1 _5042_ (.A_N(_0411_),
    .B(_0408_),
    .C(_0409_),
    .X(_0446_));
 sky130_fd_sc_hd__nand3_2 _5043_ (.A(_0403_),
    .B(_0404_),
    .C(_0405_),
    .Y(_0447_));
 sky130_fd_sc_hd__nor3_1 _5044_ (.A(_0331_),
    .B(_0400_),
    .C(_0402_),
    .Y(_0448_));
 sky130_fd_sc_hd__or2_1 _5045_ (.A(_0354_),
    .B(_0356_),
    .X(_0449_));
 sky130_fd_sc_hd__and3_1 _5046_ (.A(_1384_),
    .B(_0328_),
    .C(_0323_),
    .X(_0450_));
 sky130_fd_sc_hd__or2_1 _5047_ (.A(_0341_),
    .B(_0343_),
    .X(_0451_));
 sky130_fd_sc_hd__buf_2 _5048_ (.A(net40),
    .X(_0452_));
 sky130_fd_sc_hd__clkbuf_4 _5049_ (.A(_0452_),
    .X(_0453_));
 sky130_fd_sc_hd__clkbuf_4 _5050_ (.A(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__a22o_1 _5051_ (.A1(_0445_),
    .A2(_0327_),
    .B1(_0454_),
    .B2(_0477_),
    .X(_0456_));
 sky130_fd_sc_hd__nand4_1 _5052_ (.A(_0445_),
    .B(_0991_),
    .C(_0327_),
    .D(_0454_),
    .Y(_0457_));
 sky130_fd_sc_hd__and3_2 _5053_ (.A(_0451_),
    .B(_0456_),
    .C(_0457_),
    .X(_0458_));
 sky130_fd_sc_hd__a21oi_1 _5054_ (.A1(_0456_),
    .A2(_0457_),
    .B1(_0451_),
    .Y(_0459_));
 sky130_fd_sc_hd__nor2_1 _5055_ (.A(_0458_),
    .B(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__nand2_1 _5056_ (.A(_0450_),
    .B(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__or2_1 _5057_ (.A(_0450_),
    .B(_0460_),
    .X(_0462_));
 sky130_fd_sc_hd__nand2_1 _5058_ (.A(_0461_),
    .B(_0462_),
    .Y(_0463_));
 sky130_fd_sc_hd__xnor2_1 _5059_ (.A(_0449_),
    .B(_0463_),
    .Y(_0464_));
 sky130_fd_sc_hd__or2b_1 _5060_ (.A(_0351_),
    .B_N(_0350_),
    .X(_0465_));
 sky130_fd_sc_hd__or2b_1 _5061_ (.A(_0344_),
    .B_N(_0352_),
    .X(_0467_));
 sky130_fd_sc_hd__a21bo_1 _5062_ (.A1(_0360_),
    .A2(_0367_),
    .B1_N(_0366_),
    .X(_0468_));
 sky130_fd_sc_hd__a22oi_1 _5063_ (.A1(_3440_),
    .A2(_0339_),
    .B1(_0099_),
    .B2(_1275_),
    .Y(_0469_));
 sky130_fd_sc_hd__and4_1 _5064_ (.A(_3440_),
    .B(_0194_),
    .C(_0339_),
    .D(_0340_),
    .X(_0470_));
 sky130_fd_sc_hd__nor2_1 _5065_ (.A(_0469_),
    .B(_0470_),
    .Y(_0471_));
 sky130_fd_sc_hd__nand2_1 _5066_ (.A(_0346_),
    .B(_0219_),
    .Y(_0472_));
 sky130_fd_sc_hd__xnor2_2 _5067_ (.A(_0471_),
    .B(_0472_),
    .Y(_0473_));
 sky130_fd_sc_hd__a22o_1 _5068_ (.A1(_2423_),
    .A2(_3422_),
    .B1(_3511_),
    .B2(_2368_),
    .X(_0474_));
 sky130_fd_sc_hd__nand4_2 _5069_ (.A(_3442_),
    .B(_2434_),
    .C(_0104_),
    .D(_3511_),
    .Y(_0475_));
 sky130_fd_sc_hd__nand4_2 _5070_ (.A(_2313_),
    .B(_3619_),
    .C(_0474_),
    .D(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__a22o_1 _5071_ (.A1(_2324_),
    .A2(_0110_),
    .B1(_0474_),
    .B2(_0475_),
    .X(_0478_));
 sky130_fd_sc_hd__a32o_1 _5072_ (.A1(_0095_),
    .A2(_0110_),
    .A3(_0348_),
    .B1(_0347_),
    .B2(_3423_),
    .X(_0479_));
 sky130_fd_sc_hd__nand3_4 _5073_ (.A(_0476_),
    .B(_0478_),
    .C(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__a21o_1 _5074_ (.A1(_0476_),
    .A2(_0478_),
    .B1(_0479_),
    .X(_0481_));
 sky130_fd_sc_hd__nand3_2 _5075_ (.A(_0473_),
    .B(_0480_),
    .C(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__a21o_1 _5076_ (.A1(_0480_),
    .A2(_0481_),
    .B1(_0473_),
    .X(_0483_));
 sky130_fd_sc_hd__and3_1 _5077_ (.A(_0468_),
    .B(_0482_),
    .C(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__a21oi_1 _5078_ (.A1(_0482_),
    .A2(_0483_),
    .B1(_0468_),
    .Y(_0485_));
 sky130_fd_sc_hd__a211oi_2 _5079_ (.A1(_0465_),
    .A2(_0467_),
    .B1(_0484_),
    .C1(_0485_),
    .Y(_0486_));
 sky130_fd_sc_hd__o211a_1 _5080_ (.A1(_0484_),
    .A2(_0485_),
    .B1(_0465_),
    .C1(_0467_),
    .X(_0487_));
 sky130_fd_sc_hd__nand3_1 _5081_ (.A(_0371_),
    .B(_0392_),
    .C(_0393_),
    .Y(_0489_));
 sky130_fd_sc_hd__nand2_1 _5082_ (.A(_0363_),
    .B(_0364_),
    .Y(_0490_));
 sky130_fd_sc_hd__clkbuf_4 _5083_ (.A(net4),
    .X(_0491_));
 sky130_fd_sc_hd__a32oi_2 _5084_ (.A1(net60),
    .A2(_2204_),
    .A3(_0375_),
    .B1(_0374_),
    .B2(_0491_),
    .Y(_0492_));
 sky130_fd_sc_hd__a22o_1 _5085_ (.A1(net162),
    .A2(net32),
    .B1(net2),
    .B2(net61),
    .X(_0493_));
 sky130_fd_sc_hd__nand4_2 _5086_ (.A(_3433_),
    .B(_3431_),
    .C(net32),
    .D(net2),
    .Y(_0494_));
 sky130_fd_sc_hd__and3_1 _5087_ (.A(_3388_),
    .B(_0493_),
    .C(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__a21oi_1 _5088_ (.A1(_0493_),
    .A2(_0494_),
    .B1(_3388_),
    .Y(_0496_));
 sky130_fd_sc_hd__or3_2 _5089_ (.A(_0492_),
    .B(_0495_),
    .C(_0496_),
    .X(_0497_));
 sky130_fd_sc_hd__o21ai_1 _5090_ (.A1(_0495_),
    .A2(_0496_),
    .B1(_0492_),
    .Y(_0498_));
 sky130_fd_sc_hd__and2_1 _5091_ (.A(_0497_),
    .B(_0498_),
    .X(_0500_));
 sky130_fd_sc_hd__xor2_2 _5092_ (.A(_0490_),
    .B(_0500_),
    .X(_0501_));
 sky130_fd_sc_hd__nand2_1 _5093_ (.A(_0042_),
    .B(_2259_),
    .Y(_0502_));
 sky130_fd_sc_hd__a22oi_2 _5094_ (.A1(_0041_),
    .A2(_0491_),
    .B1(_2696_),
    .B2(_3645_),
    .Y(_0503_));
 sky130_fd_sc_hd__and4_1 _5095_ (.A(_3645_),
    .B(_0041_),
    .C(_0491_),
    .D(_2686_),
    .X(_0504_));
 sky130_fd_sc_hd__nor2_1 _5096_ (.A(_0503_),
    .B(_0504_),
    .Y(_0505_));
 sky130_fd_sc_hd__xnor2_2 _5097_ (.A(_0502_),
    .B(_0505_),
    .Y(_0506_));
 sky130_fd_sc_hd__and2_1 _5098_ (.A(_0292_),
    .B(_2740_),
    .X(_0507_));
 sky130_fd_sc_hd__a22o_1 _5099_ (.A1(_3448_),
    .A2(_0380_),
    .B1(_2489_),
    .B2(_3449_),
    .X(_0508_));
 sky130_fd_sc_hd__nand4_1 _5100_ (.A(_3451_),
    .B(_3452_),
    .C(_0380_),
    .D(_2489_),
    .Y(_0509_));
 sky130_fd_sc_hd__nand3_1 _5101_ (.A(_0507_),
    .B(_0508_),
    .C(_0509_),
    .Y(_0511_));
 sky130_fd_sc_hd__a21o_1 _5102_ (.A1(_0508_),
    .A2(_0509_),
    .B1(_0507_),
    .X(_0512_));
 sky130_fd_sc_hd__a21bo_1 _5103_ (.A1(_0378_),
    .A2(_0381_),
    .B1_N(_0382_),
    .X(_0513_));
 sky130_fd_sc_hd__nand3_2 _5104_ (.A(_0511_),
    .B(_0512_),
    .C(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__a21o_1 _5105_ (.A1(_0511_),
    .A2(_0512_),
    .B1(_0513_),
    .X(_0515_));
 sky130_fd_sc_hd__nand3_2 _5106_ (.A(_0506_),
    .B(_0514_),
    .C(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__a21o_1 _5107_ (.A1(_0514_),
    .A2(_0515_),
    .B1(_0506_),
    .X(_0517_));
 sky130_fd_sc_hd__a21bo_1 _5108_ (.A1(_0377_),
    .A2(_0387_),
    .B1_N(_0386_),
    .X(_0518_));
 sky130_fd_sc_hd__nand3_4 _5109_ (.A(_0516_),
    .B(_0517_),
    .C(_0518_),
    .Y(_0519_));
 sky130_fd_sc_hd__a21o_1 _5110_ (.A1(_0516_),
    .A2(_0517_),
    .B1(_0518_),
    .X(_0520_));
 sky130_fd_sc_hd__and3_1 _5111_ (.A(_0501_),
    .B(_0519_),
    .C(_0520_),
    .X(_0522_));
 sky130_fd_sc_hd__a21oi_1 _5112_ (.A1(_0519_),
    .A2(_0520_),
    .B1(_0501_),
    .Y(_0523_));
 sky130_fd_sc_hd__a211o_1 _5113_ (.A1(_0392_),
    .A2(_0489_),
    .B1(_0522_),
    .C1(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__o211ai_2 _5114_ (.A1(_0522_),
    .A2(_0523_),
    .B1(_0392_),
    .C1(_0489_),
    .Y(_0525_));
 sky130_fd_sc_hd__or4bb_2 _5115_ (.A(_0486_),
    .B(_0487_),
    .C_N(_0524_),
    .D_N(_0525_),
    .X(_0526_));
 sky130_fd_sc_hd__a2bb2o_1 _5116_ (.A1_N(_0486_),
    .A2_N(_0487_),
    .B1(_0524_),
    .B2(_0525_),
    .X(_0527_));
 sky130_fd_sc_hd__o211ai_4 _5117_ (.A1(net173),
    .A2(net114),
    .B1(net125),
    .C1(_0527_),
    .Y(_0528_));
 sky130_fd_sc_hd__a211o_1 _5118_ (.A1(_0526_),
    .A2(_0527_),
    .B1(net173),
    .C1(net202),
    .X(_0529_));
 sky130_fd_sc_hd__nand3_2 _5119_ (.A(_0464_),
    .B(_0528_),
    .C(_0529_),
    .Y(_0530_));
 sky130_fd_sc_hd__a21o_1 _5120_ (.A1(_0528_),
    .A2(_0529_),
    .B1(_0464_),
    .X(_0531_));
 sky130_fd_sc_hd__o211a_2 _5121_ (.A1(_0400_),
    .A2(_0448_),
    .B1(_0530_),
    .C1(_0531_),
    .X(_0533_));
 sky130_fd_sc_hd__a211oi_2 _5122_ (.A1(_0530_),
    .A2(_0531_),
    .B1(_0400_),
    .C1(_0448_),
    .Y(_0534_));
 sky130_fd_sc_hd__and2_1 _5123_ (.A(_0322_),
    .B(_0330_),
    .X(_0535_));
 sky130_fd_sc_hd__nor3b_4 _5124_ (.A(_0533_),
    .B(_0534_),
    .C_N(_0535_),
    .Y(_0536_));
 sky130_fd_sc_hd__o21ba_1 _5125_ (.A1(_0533_),
    .A2(_0534_),
    .B1_N(_0535_),
    .X(_0537_));
 sky130_fd_sc_hd__a211o_1 _5126_ (.A1(_0447_),
    .A2(_0408_),
    .B1(_0536_),
    .C1(_0537_),
    .X(_0538_));
 sky130_fd_sc_hd__o211ai_2 _5127_ (.A1(_0536_),
    .A2(_0537_),
    .B1(_0447_),
    .C1(_0408_),
    .Y(_0539_));
 sky130_fd_sc_hd__nand3_1 _5128_ (.A(_0446_),
    .B(_0538_),
    .C(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__a21o_1 _5129_ (.A1(_0538_),
    .A2(_0539_),
    .B1(_0446_),
    .X(_0541_));
 sky130_fd_sc_hd__nor3_1 _5130_ (.A(_0283_),
    .B(_0282_),
    .C(_0410_),
    .Y(_0542_));
 sky130_fd_sc_hd__and3_1 _5131_ (.A(_0540_),
    .B(_0541_),
    .C(_0542_),
    .X(_0544_));
 sky130_fd_sc_hd__a21oi_1 _5132_ (.A1(_0540_),
    .A2(_0541_),
    .B1(_0542_),
    .Y(_0545_));
 sky130_fd_sc_hd__or2_1 _5133_ (.A(_0544_),
    .B(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__or2_1 _5134_ (.A(_0321_),
    .B(_0414_),
    .X(_0547_));
 sky130_fd_sc_hd__and2_1 _5135_ (.A(_0321_),
    .B(_0414_),
    .X(_0548_));
 sky130_fd_sc_hd__a21oi_2 _5136_ (.A1(_0416_),
    .A2(_0547_),
    .B1(_0548_),
    .Y(_0549_));
 sky130_fd_sc_hd__inv_2 _5137_ (.A(_0081_),
    .Y(_0550_));
 sky130_fd_sc_hd__or2_1 _5138_ (.A(_0286_),
    .B(_0415_),
    .X(_0551_));
 sky130_fd_sc_hd__or4bb_2 _5139_ (.A(_0550_),
    .B(_0551_),
    .C_N(_0083_),
    .D_N(_0170_),
    .X(_0552_));
 sky130_fd_sc_hd__or2_1 _5140_ (.A(_0288_),
    .B(_0551_),
    .X(_0553_));
 sky130_fd_sc_hd__and3_1 _5141_ (.A(_0549_),
    .B(_0552_),
    .C(_0553_),
    .X(_0555_));
 sky130_fd_sc_hd__nand2_1 _5142_ (.A(_0546_),
    .B(_0555_),
    .Y(_0556_));
 sky130_fd_sc_hd__or2_1 _5143_ (.A(_0546_),
    .B(_0555_),
    .X(_0557_));
 sky130_fd_sc_hd__clkbuf_4 _5144_ (.A(_2510_),
    .X(_0558_));
 sky130_fd_sc_hd__clkbuf_4 _5145_ (.A(_0454_),
    .X(_0559_));
 sky130_fd_sc_hd__nor2_1 _5146_ (.A(_0558_),
    .B(_0559_),
    .Y(_0560_));
 sky130_fd_sc_hd__and2_1 _5147_ (.A(_0558_),
    .B(_0559_),
    .X(_0561_));
 sky130_fd_sc_hd__or2_1 _5148_ (.A(_0560_),
    .B(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__clkbuf_2 _5149_ (.A(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__and2b_1 _5150_ (.A_N(_0328_),
    .B(_3135_),
    .X(_0564_));
 sky130_fd_sc_hd__a31o_1 _5151_ (.A1(_3134_),
    .A2(_0337_),
    .A3(_0422_),
    .B1(_0564_),
    .X(_0566_));
 sky130_fd_sc_hd__a31o_1 _5152_ (.A1(_0296_),
    .A2(_0298_),
    .A3(_0422_),
    .B1(_0566_),
    .X(_0567_));
 sky130_fd_sc_hd__xor2_1 _5153_ (.A(_0563_),
    .B(_0567_),
    .X(_0568_));
 sky130_fd_sc_hd__nand3_1 _5154_ (.A(_0439_),
    .B(_0425_),
    .C(_0563_),
    .Y(_0569_));
 sky130_fd_sc_hd__a21o_1 _5155_ (.A1(_0439_),
    .A2(_0425_),
    .B1(_0563_),
    .X(_0570_));
 sky130_fd_sc_hd__buf_2 _5156_ (.A(net25),
    .X(_0571_));
 sky130_fd_sc_hd__mux2_1 _5157_ (.A0(_3401_),
    .A1(_3403_),
    .S(_0199_),
    .X(_0572_));
 sky130_fd_sc_hd__clkbuf_4 _5158_ (.A(_0838_),
    .X(_0573_));
 sky130_fd_sc_hd__mux2_1 _5159_ (.A0(_0571_),
    .A1(_0572_),
    .S(_0573_),
    .X(_0574_));
 sky130_fd_sc_hd__nor2_2 _5160_ (.A(_0630_),
    .B(_3154_),
    .Y(_0575_));
 sky130_fd_sc_hd__a32o_1 _5161_ (.A1(_0419_),
    .A2(_0569_),
    .A3(_0570_),
    .B1(_0574_),
    .B2(_0575_),
    .X(_0577_));
 sky130_fd_sc_hd__nor2_2 _5162_ (.A(_0783_),
    .B(_3156_),
    .Y(_0578_));
 sky130_fd_sc_hd__nand2_1 _5163_ (.A(_0558_),
    .B(_0559_),
    .Y(_0579_));
 sky130_fd_sc_hd__a21oi_1 _5164_ (.A1(_0438_),
    .A2(_0579_),
    .B1(_0000_),
    .Y(_0580_));
 sky130_fd_sc_hd__nor2_1 _5165_ (.A(_0560_),
    .B(_0580_),
    .Y(_0581_));
 sky130_fd_sc_hd__a221o_1 _5166_ (.A1(_3414_),
    .A2(_0560_),
    .B1(_0561_),
    .B2(_3194_),
    .C1(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__clkbuf_4 _5167_ (.A(_3046_),
    .X(_0583_));
 sky130_fd_sc_hd__clkbuf_4 _5168_ (.A(_3591_),
    .X(_0584_));
 sky130_fd_sc_hd__mux4_1 _5169_ (.A0(_0558_),
    .A1(_3135_),
    .A2(_3134_),
    .A3(_3133_),
    .S0(_0583_),
    .S1(_0584_),
    .X(_0585_));
 sky130_fd_sc_hd__mux4_1 _5170_ (.A0(_1078_),
    .A1(_3407_),
    .A2(_0004_),
    .A3(_0585_),
    .S0(_0429_),
    .S1(_0189_),
    .X(_0586_));
 sky130_fd_sc_hd__o21ai_1 _5171_ (.A1(_3210_),
    .A2(_0196_),
    .B1(_3727_),
    .Y(_0588_));
 sky130_fd_sc_hd__o211a_1 _5172_ (.A1(_0428_),
    .A2(_0586_),
    .B1(_0588_),
    .C1(_0849_),
    .X(_0589_));
 sky130_fd_sc_hd__a211o_1 _5173_ (.A1(_0572_),
    .A2(_0578_),
    .B1(_0582_),
    .C1(_0589_),
    .X(_0590_));
 sky130_fd_sc_hd__a211o_1 _5174_ (.A1(_3571_),
    .A2(_0568_),
    .B1(_0577_),
    .C1(_0590_),
    .X(_0591_));
 sky130_fd_sc_hd__a31o_2 _5175_ (.A1(_0320_),
    .A2(_0556_),
    .A3(_0557_),
    .B1(_0591_),
    .X(net76));
 sky130_fd_sc_hd__nand3_1 _5176_ (.A(_0540_),
    .B(_0541_),
    .C(_0542_),
    .Y(_0592_));
 sky130_fd_sc_hd__nand2_1 _5177_ (.A(_0490_),
    .B(_0500_),
    .Y(_0593_));
 sky130_fd_sc_hd__nand2_1 _5178_ (.A(_0215_),
    .B(_0219_),
    .Y(_0594_));
 sky130_fd_sc_hd__and3_1 _5179_ (.A(_3440_),
    .B(_3635_),
    .C(_0340_),
    .X(_0595_));
 sky130_fd_sc_hd__a22o_1 _5180_ (.A1(_3635_),
    .A2(net36),
    .B1(_0340_),
    .B2(_3440_),
    .X(_0596_));
 sky130_fd_sc_hd__a21bo_1 _5181_ (.A1(_3719_),
    .A2(_0595_),
    .B1_N(_0596_),
    .X(_0598_));
 sky130_fd_sc_hd__xor2_2 _5182_ (.A(_0594_),
    .B(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__a22oi_1 _5183_ (.A1(_2106_),
    .A2(_3422_),
    .B1(_0105_),
    .B2(_2434_),
    .Y(_0600_));
 sky130_fd_sc_hd__and4_1 _5184_ (.A(_2423_),
    .B(net31),
    .C(net64),
    .D(_3572_),
    .X(_0601_));
 sky130_fd_sc_hd__and4bb_1 _5185_ (.A_N(_0600_),
    .B_N(_0601_),
    .C(_2379_),
    .D(_3619_),
    .X(_0602_));
 sky130_fd_sc_hd__o2bb2a_1 _5186_ (.A1_N(_2379_),
    .A2_N(_0110_),
    .B1(_0600_),
    .B2(_0601_),
    .X(_0603_));
 sky130_fd_sc_hd__nor2_1 _5187_ (.A(_0602_),
    .B(_0603_),
    .Y(_0604_));
 sky130_fd_sc_hd__and2_1 _5188_ (.A(_0475_),
    .B(_0476_),
    .X(_0605_));
 sky130_fd_sc_hd__xnor2_2 _5189_ (.A(_0604_),
    .B(_0605_),
    .Y(_0606_));
 sky130_fd_sc_hd__xnor2_2 _5190_ (.A(_0599_),
    .B(_0606_),
    .Y(_0607_));
 sky130_fd_sc_hd__a21oi_4 _5191_ (.A1(_0497_),
    .A2(_0593_),
    .B1(_0607_),
    .Y(_0609_));
 sky130_fd_sc_hd__and3_1 _5192_ (.A(_0497_),
    .B(_0593_),
    .C(_0607_),
    .X(_0610_));
 sky130_fd_sc_hd__a211oi_4 _5193_ (.A1(_0480_),
    .A2(_0482_),
    .B1(_0609_),
    .C1(_0610_),
    .Y(_0611_));
 sky130_fd_sc_hd__o211a_1 _5194_ (.A1(_0609_),
    .A2(_0610_),
    .B1(_0480_),
    .C1(_0482_),
    .X(_0612_));
 sky130_fd_sc_hd__nand3_2 _5195_ (.A(_0501_),
    .B(_0519_),
    .C(_0520_),
    .Y(_0613_));
 sky130_fd_sc_hd__a21boi_2 _5196_ (.A1(_3388_),
    .A2(_0493_),
    .B1_N(_0494_),
    .Y(_0614_));
 sky130_fd_sc_hd__o21ba_1 _5197_ (.A1(_0502_),
    .A2(_0503_),
    .B1_N(_0504_),
    .X(_0615_));
 sky130_fd_sc_hd__a22oi_1 _5198_ (.A1(_3271_),
    .A2(_2204_),
    .B1(_2248_),
    .B2(_3632_),
    .Y(_0616_));
 sky130_fd_sc_hd__and4_1 _5199_ (.A(_3632_),
    .B(_3633_),
    .C(_3537_),
    .D(_3651_),
    .X(_0617_));
 sky130_fd_sc_hd__and4bb_1 _5200_ (.A_N(_0616_),
    .B_N(_0617_),
    .C(_3631_),
    .D(_0247_),
    .X(_0618_));
 sky130_fd_sc_hd__o2bb2a_1 _5201_ (.A1_N(_3631_),
    .A2_N(_0247_),
    .B1(_0616_),
    .B2(_0617_),
    .X(_0620_));
 sky130_fd_sc_hd__nor2_1 _5202_ (.A(_0618_),
    .B(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__xnor2_2 _5203_ (.A(_0615_),
    .B(_0621_),
    .Y(_0622_));
 sky130_fd_sc_hd__xnor2_2 _5204_ (.A(_0614_),
    .B(_0622_),
    .Y(_0623_));
 sky130_fd_sc_hd__nand2_1 _5205_ (.A(_0042_),
    .B(_2653_),
    .Y(_0624_));
 sky130_fd_sc_hd__a22oi_2 _5206_ (.A1(_0041_),
    .A2(_2696_),
    .B1(_2740_),
    .B2(_0172_),
    .Y(_0625_));
 sky130_fd_sc_hd__and4_1 _5207_ (.A(_3645_),
    .B(_0041_),
    .C(_2686_),
    .D(_2740_),
    .X(_0626_));
 sky130_fd_sc_hd__nor2_1 _5208_ (.A(_0625_),
    .B(_0626_),
    .Y(_0627_));
 sky130_fd_sc_hd__xnor2_2 _5209_ (.A(_0624_),
    .B(_0627_),
    .Y(_0628_));
 sky130_fd_sc_hd__and2_1 _5210_ (.A(_0292_),
    .B(_0380_),
    .X(_0629_));
 sky130_fd_sc_hd__a22o_1 _5211_ (.A1(_3452_),
    .A2(_2489_),
    .B1(_2521_),
    .B2(_3449_),
    .X(_0631_));
 sky130_fd_sc_hd__nand4_1 _5212_ (.A(_3451_),
    .B(_3452_),
    .C(_2489_),
    .D(_2521_),
    .Y(_0632_));
 sky130_fd_sc_hd__nand3_1 _5213_ (.A(_0629_),
    .B(_0631_),
    .C(_0632_),
    .Y(_0633_));
 sky130_fd_sc_hd__a21o_1 _5214_ (.A1(_0631_),
    .A2(_0632_),
    .B1(_0629_),
    .X(_0634_));
 sky130_fd_sc_hd__a21bo_1 _5215_ (.A1(_0507_),
    .A2(_0508_),
    .B1_N(_0509_),
    .X(_0635_));
 sky130_fd_sc_hd__nand3_2 _5216_ (.A(_0633_),
    .B(_0634_),
    .C(_0635_),
    .Y(_0636_));
 sky130_fd_sc_hd__a21o_1 _5217_ (.A1(_0633_),
    .A2(_0634_),
    .B1(_0635_),
    .X(_0637_));
 sky130_fd_sc_hd__nand3_2 _5218_ (.A(_0628_),
    .B(_0636_),
    .C(_0637_),
    .Y(_0638_));
 sky130_fd_sc_hd__a21o_1 _5219_ (.A1(_0636_),
    .A2(_0637_),
    .B1(_0628_),
    .X(_0639_));
 sky130_fd_sc_hd__a21bo_1 _5220_ (.A1(_0506_),
    .A2(_0515_),
    .B1_N(_0514_),
    .X(_0640_));
 sky130_fd_sc_hd__nand3_4 _5221_ (.A(_0638_),
    .B(_0639_),
    .C(_0640_),
    .Y(_0642_));
 sky130_fd_sc_hd__a21o_1 _5222_ (.A1(_0638_),
    .A2(_0639_),
    .B1(_0640_),
    .X(_0643_));
 sky130_fd_sc_hd__and3_1 _5223_ (.A(_0623_),
    .B(_0642_),
    .C(_0643_),
    .X(_0644_));
 sky130_fd_sc_hd__a21oi_2 _5224_ (.A1(_0642_),
    .A2(_0643_),
    .B1(_0623_),
    .Y(_0645_));
 sky130_fd_sc_hd__a211oi_4 _5225_ (.A1(_0519_),
    .A2(_0613_),
    .B1(_0644_),
    .C1(_0645_),
    .Y(_0646_));
 sky130_fd_sc_hd__o211a_1 _5226_ (.A1(_0644_),
    .A2(_0645_),
    .B1(_0519_),
    .C1(_0613_),
    .X(_0647_));
 sky130_fd_sc_hd__nor4_1 _5227_ (.A(_0611_),
    .B(_0612_),
    .C(_0646_),
    .D(_0647_),
    .Y(_0648_));
 sky130_fd_sc_hd__o22a_1 _5228_ (.A1(_0611_),
    .A2(_0612_),
    .B1(_0646_),
    .B2(_0647_),
    .X(_0649_));
 sky130_fd_sc_hd__a211oi_2 _5229_ (.A1(_0524_),
    .A2(_0526_),
    .B1(net113),
    .C1(_0649_),
    .Y(_0650_));
 sky130_fd_sc_hd__o211a_1 _5230_ (.A1(_0648_),
    .A2(_0649_),
    .B1(_0524_),
    .C1(_0526_),
    .X(_0651_));
 sky130_fd_sc_hd__and3_1 _5231_ (.A(_0346_),
    .B(_0220_),
    .C(_0471_),
    .X(_0653_));
 sky130_fd_sc_hd__buf_2 _5232_ (.A(net41),
    .X(_0654_));
 sky130_fd_sc_hd__nand2_1 _5233_ (.A(_0466_),
    .B(_0654_),
    .Y(_0655_));
 sky130_fd_sc_hd__and3_1 _5234_ (.A(_0324_),
    .B(net163),
    .C(_0452_),
    .X(_0656_));
 sky130_fd_sc_hd__a22o_1 _5235_ (.A1(_0324_),
    .A2(_0325_),
    .B1(_0453_),
    .B2(net163),
    .X(_0657_));
 sky130_fd_sc_hd__a21bo_1 _5236_ (.A1(_0326_),
    .A2(_0656_),
    .B1_N(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__xor2_1 _5237_ (.A(_0655_),
    .B(_0658_),
    .X(_0659_));
 sky130_fd_sc_hd__o21a_1 _5238_ (.A1(_0470_),
    .A2(_0653_),
    .B1(_0659_),
    .X(_0660_));
 sky130_fd_sc_hd__or3_1 _5239_ (.A(_0470_),
    .B(_0653_),
    .C(_0659_),
    .X(_0661_));
 sky130_fd_sc_hd__and2b_1 _5240_ (.A_N(_0660_),
    .B(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__and4_1 _5241_ (.A(_0445_),
    .B(_0991_),
    .C(_0327_),
    .D(_0454_),
    .X(_0664_));
 sky130_fd_sc_hd__nor2_1 _5242_ (.A(_0664_),
    .B(_0458_),
    .Y(_0665_));
 sky130_fd_sc_hd__xnor2_1 _5243_ (.A(_0662_),
    .B(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__o21ai_1 _5244_ (.A1(_0484_),
    .A2(_0486_),
    .B1(_0666_),
    .Y(_0667_));
 sky130_fd_sc_hd__or3_1 _5245_ (.A(_0484_),
    .B(_0486_),
    .C(_0666_),
    .X(_0668_));
 sky130_fd_sc_hd__nand2_1 _5246_ (.A(_0667_),
    .B(_0668_),
    .Y(_0669_));
 sky130_fd_sc_hd__xor2_1 _5247_ (.A(_0461_),
    .B(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__nor3b_2 _5248_ (.A(_0650_),
    .B(_0651_),
    .C_N(_0670_),
    .Y(_0671_));
 sky130_fd_sc_hd__o21ba_1 _5249_ (.A1(_0650_),
    .A2(_0651_),
    .B1_N(_0670_),
    .X(_0672_));
 sky130_fd_sc_hd__a211oi_2 _5250_ (.A1(_0528_),
    .A2(_0530_),
    .B1(_0671_),
    .C1(_0672_),
    .Y(_0673_));
 sky130_fd_sc_hd__o211a_1 _5251_ (.A1(_0671_),
    .A2(_0672_),
    .B1(_0528_),
    .C1(_0530_),
    .X(_0675_));
 sky130_fd_sc_hd__and2b_1 _5252_ (.A_N(_0463_),
    .B(_0449_),
    .X(_0676_));
 sky130_fd_sc_hd__or3b_1 _5253_ (.A(_0673_),
    .B(_0675_),
    .C_N(_0676_),
    .X(_0677_));
 sky130_fd_sc_hd__o21bai_1 _5254_ (.A1(_0673_),
    .A2(_0675_),
    .B1_N(_0676_),
    .Y(_0678_));
 sky130_fd_sc_hd__o211a_1 _5255_ (.A1(_0533_),
    .A2(_0536_),
    .B1(_0677_),
    .C1(_0678_),
    .X(_0679_));
 sky130_fd_sc_hd__a211o_1 _5256_ (.A1(_0677_),
    .A2(_0678_),
    .B1(_0533_),
    .C1(_0536_),
    .X(_0680_));
 sky130_fd_sc_hd__or2b_1 _5257_ (.A(_0679_),
    .B_N(_0680_),
    .X(_0681_));
 sky130_fd_sc_hd__a211oi_2 _5258_ (.A1(_0447_),
    .A2(_0408_),
    .B1(_0536_),
    .C1(_0537_),
    .Y(_0682_));
 sky130_fd_sc_hd__a21oi_1 _5259_ (.A1(_0446_),
    .A2(_0539_),
    .B1(_0682_),
    .Y(_0683_));
 sky130_fd_sc_hd__xnor2_1 _5260_ (.A(_0681_),
    .B(_0683_),
    .Y(_0684_));
 sky130_fd_sc_hd__a21oi_1 _5261_ (.A1(_0592_),
    .A2(_0557_),
    .B1(_0684_),
    .Y(_0686_));
 sky130_fd_sc_hd__a31o_1 _5262_ (.A1(_0592_),
    .A2(_0557_),
    .A3(_0684_),
    .B1(_3192_),
    .X(_0687_));
 sky130_fd_sc_hd__clkbuf_4 _5263_ (.A(_0654_),
    .X(_0688_));
 sky130_fd_sc_hd__clkbuf_4 _5264_ (.A(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__and2_1 _5265_ (.A(_3128_),
    .B(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__nor2_1 _5266_ (.A(_3128_),
    .B(_0689_),
    .Y(_0691_));
 sky130_fd_sc_hd__or2_1 _5267_ (.A(_0690_),
    .B(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__clkbuf_2 _5268_ (.A(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__and2b_1 _5269_ (.A_N(_0559_),
    .B(_0558_),
    .X(_0694_));
 sky130_fd_sc_hd__a21o_1 _5270_ (.A1(_0563_),
    .A2(_0567_),
    .B1(_0694_),
    .X(_0695_));
 sky130_fd_sc_hd__xor2_1 _5271_ (.A(_0693_),
    .B(_0695_),
    .X(_0697_));
 sky130_fd_sc_hd__nand2_2 _5272_ (.A(_3571_),
    .B(_0697_),
    .Y(_0698_));
 sky130_fd_sc_hd__a21oi_1 _5273_ (.A1(_0579_),
    .A2(_0570_),
    .B1(_0693_),
    .Y(_0699_));
 sky130_fd_sc_hd__a31o_1 _5274_ (.A1(_0579_),
    .A2(_0570_),
    .A3(_0693_),
    .B1(_3596_),
    .X(_0700_));
 sky130_fd_sc_hd__mux2_1 _5275_ (.A0(_3132_),
    .A1(_3151_),
    .S(_1100_),
    .X(_0701_));
 sky130_fd_sc_hd__a211o_1 _5276_ (.A1(_1100_),
    .A2(_3145_),
    .B1(_3492_),
    .C1(_1723_),
    .X(_0702_));
 sky130_fd_sc_hd__a21bo_1 _5277_ (.A1(_1723_),
    .A2(_0701_),
    .B1_N(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__or2_1 _5278_ (.A(_3128_),
    .B(_0689_),
    .X(_0704_));
 sky130_fd_sc_hd__o21bai_1 _5279_ (.A1(_3589_),
    .A2(_0690_),
    .B1_N(_0000_),
    .Y(_0705_));
 sky130_fd_sc_hd__a31o_1 _5280_ (.A1(_0583_),
    .A2(_0584_),
    .A3(_1734_),
    .B1(_3580_),
    .X(_0706_));
 sky130_fd_sc_hd__a22o_1 _5281_ (.A1(_3194_),
    .A2(_0690_),
    .B1(_0691_),
    .B2(_3414_),
    .X(_0708_));
 sky130_fd_sc_hd__a221o_1 _5282_ (.A1(_0704_),
    .A2(_0705_),
    .B1(_0706_),
    .B2(_3161_),
    .C1(_0708_),
    .X(_0709_));
 sky130_fd_sc_hd__mux4_1 _5283_ (.A0(_3128_),
    .A1(_0558_),
    .A2(_3135_),
    .A3(_3134_),
    .S0(_3046_),
    .S1(_0584_),
    .X(_0710_));
 sky130_fd_sc_hd__mux4_1 _5284_ (.A0(_3066_),
    .A1(_3500_),
    .A2(_0187_),
    .A3(_0710_),
    .S0(_0429_),
    .S1(_0189_),
    .X(_0711_));
 sky130_fd_sc_hd__or2_1 _5285_ (.A(_3056_),
    .B(_0196_),
    .X(_0712_));
 sky130_fd_sc_hd__nand2_1 _5286_ (.A(_3727_),
    .B(_0712_),
    .Y(_0713_));
 sky130_fd_sc_hd__o211a_1 _5287_ (.A1(_3727_),
    .A2(_0711_),
    .B1(_0713_),
    .C1(_0849_),
    .X(_0714_));
 sky130_fd_sc_hd__a311o_1 _5288_ (.A1(_0573_),
    .A2(_3587_),
    .A3(_0703_),
    .B1(_0709_),
    .C1(_0714_),
    .X(_0715_));
 sky130_fd_sc_hd__o21ba_2 _5289_ (.A1(_0699_),
    .A2(_0700_),
    .B1_N(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__o211ai_4 _5290_ (.A1(_0686_),
    .A2(_0687_),
    .B1(_0698_),
    .C1(_0716_),
    .Y(net77));
 sky130_fd_sc_hd__nor3b_1 _5291_ (.A(_0673_),
    .B(_0675_),
    .C_N(_0676_),
    .Y(_0718_));
 sky130_fd_sc_hd__o21a_1 _5292_ (.A1(_0461_),
    .A2(_0669_),
    .B1(_0667_),
    .X(_0719_));
 sky130_fd_sc_hd__buf_2 _5293_ (.A(net42),
    .X(_0720_));
 sky130_fd_sc_hd__buf_2 _5294_ (.A(_0720_),
    .X(_0721_));
 sky130_fd_sc_hd__clkbuf_4 _5295_ (.A(_0721_),
    .X(_0722_));
 sky130_fd_sc_hd__nand2_2 _5296_ (.A(_1002_),
    .B(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__a32o_1 _5297_ (.A1(_0477_),
    .A2(_0688_),
    .A3(_0657_),
    .B1(_0656_),
    .B2(_0327_),
    .X(_0724_));
 sky130_fd_sc_hd__a32oi_2 _5298_ (.A1(_0205_),
    .A2(net38),
    .A3(_0596_),
    .B1(_0595_),
    .B2(_3718_),
    .Y(_0725_));
 sky130_fd_sc_hd__a22oi_1 _5299_ (.A1(_0194_),
    .A2(_0325_),
    .B1(_0452_),
    .B2(_0324_),
    .Y(_0726_));
 sky130_fd_sc_hd__and4_1 _5300_ (.A(_0194_),
    .B(_0324_),
    .C(_0325_),
    .D(_0452_),
    .X(_0727_));
 sky130_fd_sc_hd__and4bb_1 _5301_ (.A_N(_0726_),
    .B_N(_0727_),
    .C(_0423_),
    .D(net41),
    .X(_0729_));
 sky130_fd_sc_hd__o2bb2a_1 _5302_ (.A1_N(_0423_),
    .A2_N(_0654_),
    .B1(_0726_),
    .B2(_0727_),
    .X(_0730_));
 sky130_fd_sc_hd__or3_1 _5303_ (.A(_0725_),
    .B(_0729_),
    .C(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__o21ai_1 _5304_ (.A1(_0729_),
    .A2(_0730_),
    .B1(_0725_),
    .Y(_0732_));
 sky130_fd_sc_hd__and2_1 _5305_ (.A(_0731_),
    .B(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__xor2_2 _5306_ (.A(_0724_),
    .B(_0733_),
    .X(_0734_));
 sky130_fd_sc_hd__o21a_1 _5307_ (.A1(_0664_),
    .A2(_0660_),
    .B1(_0661_),
    .X(_0735_));
 sky130_fd_sc_hd__xnor2_1 _5308_ (.A(_0734_),
    .B(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__xor2_1 _5309_ (.A(_0723_),
    .B(_0736_),
    .X(_0737_));
 sky130_fd_sc_hd__o21ai_2 _5310_ (.A1(_0609_),
    .A2(_0611_),
    .B1(_0737_),
    .Y(_0738_));
 sky130_fd_sc_hd__or3_1 _5311_ (.A(_0609_),
    .B(_0611_),
    .C(_0737_),
    .X(_0740_));
 sky130_fd_sc_hd__a22o_1 _5312_ (.A1(_0458_),
    .A2(_0662_),
    .B1(_0738_),
    .B2(_0740_),
    .X(_0741_));
 sky130_fd_sc_hd__nand4_2 _5313_ (.A(_0458_),
    .B(_0662_),
    .C(_0738_),
    .D(_0740_),
    .Y(_0742_));
 sky130_fd_sc_hd__inv_2 _5314_ (.A(_0646_),
    .Y(_0743_));
 sky130_fd_sc_hd__or4_1 _5315_ (.A(_0611_),
    .B(_0612_),
    .C(_0646_),
    .D(_0647_),
    .X(_0744_));
 sky130_fd_sc_hd__and2b_1 _5316_ (.A_N(_0605_),
    .B(_0604_),
    .X(_0745_));
 sky130_fd_sc_hd__and2_1 _5317_ (.A(_0599_),
    .B(_0606_),
    .X(_0746_));
 sky130_fd_sc_hd__or3_1 _5318_ (.A(_0615_),
    .B(_0618_),
    .C(_0620_),
    .X(_0747_));
 sky130_fd_sc_hd__or2b_1 _5319_ (.A(_0614_),
    .B_N(_0622_),
    .X(_0748_));
 sky130_fd_sc_hd__a22o_1 _5320_ (.A1(_3442_),
    .A2(net36),
    .B1(net37),
    .B2(_3635_),
    .X(_0749_));
 sky130_fd_sc_hd__nand4_4 _5321_ (.A(_3635_),
    .B(_3442_),
    .C(_0339_),
    .D(_0340_),
    .Y(_0751_));
 sky130_fd_sc_hd__nand4_2 _5322_ (.A(_0095_),
    .B(net38),
    .C(_0749_),
    .D(_0751_),
    .Y(_0752_));
 sky130_fd_sc_hd__a22o_1 _5323_ (.A1(_0106_),
    .A2(_0220_),
    .B1(_0749_),
    .B2(_0751_),
    .X(_0753_));
 sky130_fd_sc_hd__and2_1 _5324_ (.A(_0752_),
    .B(_0753_),
    .X(_0754_));
 sky130_fd_sc_hd__nand2_1 _5325_ (.A(_3530_),
    .B(_0110_),
    .Y(_0755_));
 sky130_fd_sc_hd__a22oi_2 _5326_ (.A1(_0247_),
    .A2(_0104_),
    .B1(_3512_),
    .B2(_3644_),
    .Y(_0756_));
 sky130_fd_sc_hd__and4_1 _5327_ (.A(_3644_),
    .B(_2149_),
    .C(_0104_),
    .D(_0105_),
    .X(_0757_));
 sky130_fd_sc_hd__nor2_1 _5328_ (.A(_0756_),
    .B(_0757_),
    .Y(_0758_));
 sky130_fd_sc_hd__xnor2_2 _5329_ (.A(_0755_),
    .B(_0758_),
    .Y(_0759_));
 sky130_fd_sc_hd__nor2_1 _5330_ (.A(_0601_),
    .B(_0602_),
    .Y(_0760_));
 sky130_fd_sc_hd__xnor2_2 _5331_ (.A(_0759_),
    .B(_0760_),
    .Y(_0762_));
 sky130_fd_sc_hd__xnor2_2 _5332_ (.A(_0754_),
    .B(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__a21o_2 _5333_ (.A1(_0747_),
    .A2(_0748_),
    .B1(_0763_),
    .X(_0764_));
 sky130_fd_sc_hd__nand3_2 _5334_ (.A(_0747_),
    .B(_0748_),
    .C(_0763_),
    .Y(_0765_));
 sky130_fd_sc_hd__o211a_1 _5335_ (.A1(_0745_),
    .A2(_0746_),
    .B1(_0764_),
    .C1(_0765_),
    .X(_0766_));
 sky130_fd_sc_hd__a211oi_2 _5336_ (.A1(_0764_),
    .A2(_0765_),
    .B1(_0745_),
    .C1(_0746_),
    .Y(_0767_));
 sky130_fd_sc_hd__nand3_2 _5337_ (.A(_0623_),
    .B(_0642_),
    .C(_0643_),
    .Y(_0768_));
 sky130_fd_sc_hd__or2_1 _5338_ (.A(_0617_),
    .B(_0618_),
    .X(_0769_));
 sky130_fd_sc_hd__o21ba_1 _5339_ (.A1(_0624_),
    .A2(_0625_),
    .B1_N(_0626_),
    .X(_0770_));
 sky130_fd_sc_hd__a22oi_1 _5340_ (.A1(_3271_),
    .A2(_2248_),
    .B1(_0491_),
    .B2(_3196_),
    .Y(_0771_));
 sky130_fd_sc_hd__and4_1 _5341_ (.A(_3632_),
    .B(_3271_),
    .C(_3651_),
    .D(_0491_),
    .X(_0773_));
 sky130_fd_sc_hd__and4bb_1 _5342_ (.A_N(_0771_),
    .B_N(_0773_),
    .C(_3631_),
    .D(_2215_),
    .X(_0774_));
 sky130_fd_sc_hd__o2bb2a_1 _5343_ (.A1_N(_3385_),
    .A2_N(_2215_),
    .B1(_0771_),
    .B2(_0773_),
    .X(_0775_));
 sky130_fd_sc_hd__nor2_1 _5344_ (.A(_0774_),
    .B(_0775_),
    .Y(_0776_));
 sky130_fd_sc_hd__xnor2_2 _5345_ (.A(_0770_),
    .B(_0776_),
    .Y(_0777_));
 sky130_fd_sc_hd__xor2_2 _5346_ (.A(_0769_),
    .B(_0777_),
    .X(_0778_));
 sky130_fd_sc_hd__nand2_1 _5347_ (.A(_0042_),
    .B(_2696_),
    .Y(_0779_));
 sky130_fd_sc_hd__and3_1 _5348_ (.A(_0161_),
    .B(_3531_),
    .C(net6),
    .X(_0780_));
 sky130_fd_sc_hd__a22o_1 _5349_ (.A1(_3531_),
    .A2(net6),
    .B1(_0380_),
    .B2(_0161_),
    .X(_0781_));
 sky130_fd_sc_hd__a21bo_1 _5350_ (.A1(_2773_),
    .A2(_0780_),
    .B1_N(_0781_),
    .X(_0782_));
 sky130_fd_sc_hd__xor2_2 _5351_ (.A(_0779_),
    .B(_0782_),
    .X(_0784_));
 sky130_fd_sc_hd__and2_1 _5352_ (.A(_0292_),
    .B(net8),
    .X(_0785_));
 sky130_fd_sc_hd__a22o_1 _5353_ (.A1(_0390_),
    .A2(_2521_),
    .B1(net10),
    .B2(_0488_),
    .X(_0786_));
 sky130_fd_sc_hd__nand4_2 _5354_ (.A(_3449_),
    .B(_3448_),
    .C(_2521_),
    .D(_2565_),
    .Y(_0787_));
 sky130_fd_sc_hd__nand3_1 _5355_ (.A(_0785_),
    .B(_0786_),
    .C(_0787_),
    .Y(_0788_));
 sky130_fd_sc_hd__a21o_1 _5356_ (.A1(_0786_),
    .A2(_0787_),
    .B1(_0785_),
    .X(_0789_));
 sky130_fd_sc_hd__a21bo_1 _5357_ (.A1(_0629_),
    .A2(_0631_),
    .B1_N(_0632_),
    .X(_0790_));
 sky130_fd_sc_hd__nand3_1 _5358_ (.A(_0788_),
    .B(_0789_),
    .C(_0790_),
    .Y(_0791_));
 sky130_fd_sc_hd__a21o_1 _5359_ (.A1(_0788_),
    .A2(_0789_),
    .B1(_0790_),
    .X(_0792_));
 sky130_fd_sc_hd__nand3_2 _5360_ (.A(_0784_),
    .B(_0791_),
    .C(_0792_),
    .Y(_0793_));
 sky130_fd_sc_hd__a21o_1 _5361_ (.A1(_0791_),
    .A2(_0792_),
    .B1(_0784_),
    .X(_0795_));
 sky130_fd_sc_hd__a21bo_1 _5362_ (.A1(_0628_),
    .A2(_0637_),
    .B1_N(_0636_),
    .X(_0796_));
 sky130_fd_sc_hd__nand3_4 _5363_ (.A(_0793_),
    .B(_0795_),
    .C(_0796_),
    .Y(_0797_));
 sky130_fd_sc_hd__a21o_1 _5364_ (.A1(_0793_),
    .A2(_0795_),
    .B1(_0796_),
    .X(_0798_));
 sky130_fd_sc_hd__and3_1 _5365_ (.A(_0778_),
    .B(_0797_),
    .C(_0798_),
    .X(_0799_));
 sky130_fd_sc_hd__a21oi_2 _5366_ (.A1(_0797_),
    .A2(_0798_),
    .B1(_0778_),
    .Y(_0800_));
 sky130_fd_sc_hd__a211oi_4 _5367_ (.A1(_0642_),
    .A2(_0768_),
    .B1(_0799_),
    .C1(_0800_),
    .Y(_0801_));
 sky130_fd_sc_hd__o211a_1 _5368_ (.A1(_0799_),
    .A2(_0800_),
    .B1(_0642_),
    .C1(_0768_),
    .X(_0802_));
 sky130_fd_sc_hd__nor4_2 _5369_ (.A(_0766_),
    .B(_0767_),
    .C(_0801_),
    .D(_0802_),
    .Y(_0803_));
 sky130_fd_sc_hd__o22a_1 _5370_ (.A1(_0766_),
    .A2(_0767_),
    .B1(_0801_),
    .B2(_0802_),
    .X(_0804_));
 sky130_fd_sc_hd__a211o_1 _5371_ (.A1(_0743_),
    .A2(_0744_),
    .B1(net112),
    .C1(_0804_),
    .X(_0806_));
 sky130_fd_sc_hd__o211ai_2 _5372_ (.A1(net112),
    .A2(_0804_),
    .B1(_0743_),
    .C1(_0744_),
    .Y(_0807_));
 sky130_fd_sc_hd__nand4_2 _5373_ (.A(_0741_),
    .B(_0742_),
    .C(_0806_),
    .D(_0807_),
    .Y(_0808_));
 sky130_fd_sc_hd__a22o_1 _5374_ (.A1(_0741_),
    .A2(_0742_),
    .B1(_0806_),
    .B2(_0807_),
    .X(_0809_));
 sky130_fd_sc_hd__o211a_1 _5375_ (.A1(net135),
    .A2(_0671_),
    .B1(_0808_),
    .C1(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__a211oi_2 _5376_ (.A1(_0808_),
    .A2(_0809_),
    .B1(net135),
    .C1(_0671_),
    .Y(_0811_));
 sky130_fd_sc_hd__or3_1 _5377_ (.A(_0719_),
    .B(_0810_),
    .C(_0811_),
    .X(_0812_));
 sky130_fd_sc_hd__o21ai_1 _5378_ (.A1(_0810_),
    .A2(_0811_),
    .B1(_0719_),
    .Y(_0813_));
 sky130_fd_sc_hd__o211a_2 _5379_ (.A1(_0673_),
    .A2(_0718_),
    .B1(_0812_),
    .C1(_0813_),
    .X(_0814_));
 sky130_fd_sc_hd__a211o_1 _5380_ (.A1(_0812_),
    .A2(_0813_),
    .B1(_0673_),
    .C1(_0718_),
    .X(_0815_));
 sky130_fd_sc_hd__nor2b_1 _5381_ (.A(_0814_),
    .B_N(_0815_),
    .Y(_0817_));
 sky130_fd_sc_hd__a21o_1 _5382_ (.A1(_0682_),
    .A2(_0680_),
    .B1(net140),
    .X(_0818_));
 sky130_fd_sc_hd__xnor2_1 _5383_ (.A(_0817_),
    .B(_0818_),
    .Y(_0819_));
 sky130_fd_sc_hd__o22a_1 _5384_ (.A1(_0540_),
    .A2(_0681_),
    .B1(_0684_),
    .B2(_0592_),
    .X(_0820_));
 sky130_fd_sc_hd__or3_1 _5385_ (.A(_0544_),
    .B(_0545_),
    .C(_0684_),
    .X(_0821_));
 sky130_fd_sc_hd__a31o_1 _5386_ (.A1(_0549_),
    .A2(_0552_),
    .A3(_0553_),
    .B1(_0821_),
    .X(_0822_));
 sky130_fd_sc_hd__and3_1 _5387_ (.A(_0819_),
    .B(_0820_),
    .C(_0822_),
    .X(_0823_));
 sky130_fd_sc_hd__a21oi_1 _5388_ (.A1(_0820_),
    .A2(_0822_),
    .B1(_0819_),
    .Y(_0824_));
 sky130_fd_sc_hd__or2_1 _5389_ (.A(_3192_),
    .B(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__and2_2 _5390_ (.A(_2587_),
    .B(_0722_),
    .X(_0826_));
 sky130_fd_sc_hd__nor2_1 _5391_ (.A(_2587_),
    .B(_0722_),
    .Y(_0828_));
 sky130_fd_sc_hd__or2_2 _5392_ (.A(_0826_),
    .B(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__and2b_1 _5393_ (.A_N(_0689_),
    .B(_3128_),
    .X(_0830_));
 sky130_fd_sc_hd__a21o_1 _5394_ (.A1(_0693_),
    .A2(_0695_),
    .B1(_0830_),
    .X(_0831_));
 sky130_fd_sc_hd__nor2_1 _5395_ (.A(_0829_),
    .B(_0831_),
    .Y(_0832_));
 sky130_fd_sc_hd__and2_1 _5396_ (.A(_0829_),
    .B(_0831_),
    .X(_0833_));
 sky130_fd_sc_hd__a31oi_2 _5397_ (.A1(_0558_),
    .A2(_0559_),
    .A3(_0704_),
    .B1(_0690_),
    .Y(_0834_));
 sky130_fd_sc_hd__a211o_1 _5398_ (.A1(_0439_),
    .A2(_0425_),
    .B1(_0563_),
    .C1(_0693_),
    .X(_0835_));
 sky130_fd_sc_hd__a21oi_2 _5399_ (.A1(_0834_),
    .A2(_0835_),
    .B1(_0829_),
    .Y(_0836_));
 sky130_fd_sc_hd__a311o_1 _5400_ (.A1(_0829_),
    .A2(_0834_),
    .A3(_0835_),
    .B1(_0836_),
    .C1(_3596_),
    .X(_0837_));
 sky130_fd_sc_hd__mux2_1 _5401_ (.A0(_3582_),
    .A1(_3584_),
    .S(_0199_),
    .X(_0839_));
 sky130_fd_sc_hd__or2_1 _5402_ (.A(_3727_),
    .B(_3707_),
    .X(_0840_));
 sky130_fd_sc_hd__or2_1 _5403_ (.A(_0199_),
    .B(_3727_),
    .X(_0841_));
 sky130_fd_sc_hd__a32o_1 _5404_ (.A1(_0571_),
    .A2(_0840_),
    .A3(_0841_),
    .B1(_0839_),
    .B2(_0573_),
    .X(_0842_));
 sky130_fd_sc_hd__and2_1 _5405_ (.A(_0575_),
    .B(_0842_),
    .X(_0843_));
 sky130_fd_sc_hd__buf_2 _5406_ (.A(_0849_),
    .X(_0844_));
 sky130_fd_sc_hd__mux4_1 _5407_ (.A0(_2587_),
    .A1(_3128_),
    .A2(_0558_),
    .A3(_3135_),
    .S0(_0583_),
    .S1(_0584_),
    .X(_0845_));
 sky130_fd_sc_hd__mux4_1 _5408_ (.A0(_3207_),
    .A1(_3602_),
    .A2(_0304_),
    .A3(_0845_),
    .S0(_0429_),
    .S1(_0189_),
    .X(_0846_));
 sky130_fd_sc_hd__or2_1 _5409_ (.A(_0428_),
    .B(_0846_),
    .X(_0847_));
 sky130_fd_sc_hd__buf_2 _5410_ (.A(_0428_),
    .X(_0848_));
 sky130_fd_sc_hd__nand2_2 _5411_ (.A(_3212_),
    .B(_3729_),
    .Y(_0850_));
 sky130_fd_sc_hd__nand2_1 _5412_ (.A(_0848_),
    .B(_0850_),
    .Y(_0851_));
 sky130_fd_sc_hd__o21ba_1 _5413_ (.A1(_3589_),
    .A2(_0826_),
    .B1_N(_0000_),
    .X(_0852_));
 sky130_fd_sc_hd__nor2_1 _5414_ (.A(_0828_),
    .B(_0852_),
    .Y(_0853_));
 sky130_fd_sc_hd__clkbuf_4 _5415_ (.A(_3194_),
    .X(_0854_));
 sky130_fd_sc_hd__clkbuf_4 _5416_ (.A(_3414_),
    .X(_0855_));
 sky130_fd_sc_hd__a22o_1 _5417_ (.A1(_0854_),
    .A2(_0826_),
    .B1(_0828_),
    .B2(_0855_),
    .X(_0856_));
 sky130_fd_sc_hd__a311o_1 _5418_ (.A1(_0844_),
    .A2(_0847_),
    .A3(_0851_),
    .B1(_0853_),
    .C1(_0856_),
    .X(_0857_));
 sky130_fd_sc_hd__a211oi_1 _5419_ (.A1(_0578_),
    .A2(_0839_),
    .B1(_0843_),
    .C1(_0857_),
    .Y(_0858_));
 sky130_fd_sc_hd__o311a_2 _5420_ (.A1(_0181_),
    .A2(_0832_),
    .A3(_0833_),
    .B1(_0837_),
    .C1(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__o21ai_4 _5421_ (.A1(_0823_),
    .A2(_0825_),
    .B1(_0859_),
    .Y(net78));
 sky130_fd_sc_hd__clkbuf_4 _5422_ (.A(_0848_),
    .X(_0861_));
 sky130_fd_sc_hd__clkbuf_4 _5423_ (.A(_2609_),
    .X(_0862_));
 sky130_fd_sc_hd__buf_4 _5424_ (.A(_0583_),
    .X(_0863_));
 sky130_fd_sc_hd__clkbuf_4 _5425_ (.A(_0584_),
    .X(_0864_));
 sky130_fd_sc_hd__mux4_1 _5426_ (.A0(_0862_),
    .A1(_2587_),
    .A2(_3128_),
    .A3(_0558_),
    .S0(_0863_),
    .S1(_0864_),
    .X(_0865_));
 sky130_fd_sc_hd__clkbuf_4 _5427_ (.A(_0429_),
    .X(_0866_));
 sky130_fd_sc_hd__clkbuf_4 _5428_ (.A(_0189_),
    .X(_0867_));
 sky130_fd_sc_hd__mux4_1 _5429_ (.A0(_3283_),
    .A1(_3702_),
    .A2(_0433_),
    .A3(_0865_),
    .S0(_0866_),
    .S1(_0867_),
    .X(_0868_));
 sky130_fd_sc_hd__nand2_1 _5430_ (.A(_3284_),
    .B(_3729_),
    .Y(_0869_));
 sky130_fd_sc_hd__nand2_1 _5431_ (.A(_0848_),
    .B(_0869_),
    .Y(_0871_));
 sky130_fd_sc_hd__o211a_1 _5432_ (.A1(_0861_),
    .A2(_0868_),
    .B1(_0871_),
    .C1(_0844_),
    .X(_0872_));
 sky130_fd_sc_hd__buf_2 _5433_ (.A(net43),
    .X(_0873_));
 sky130_fd_sc_hd__buf_2 _5434_ (.A(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__buf_2 _5435_ (.A(_0874_),
    .X(_0875_));
 sky130_fd_sc_hd__nor2_1 _5436_ (.A(_0862_),
    .B(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__and2_2 _5437_ (.A(_0862_),
    .B(_0875_),
    .X(_0877_));
 sky130_fd_sc_hd__or2_2 _5438_ (.A(_0876_),
    .B(_0877_),
    .X(_0878_));
 sky130_fd_sc_hd__o21bai_1 _5439_ (.A1(_0826_),
    .A2(_0836_),
    .B1_N(_0878_),
    .Y(_0879_));
 sky130_fd_sc_hd__or3b_1 _5440_ (.A(_0826_),
    .B(_0836_),
    .C_N(_0878_),
    .X(_0880_));
 sky130_fd_sc_hd__mux2_1 _5441_ (.A0(_3296_),
    .A1(_3292_),
    .S(_0980_),
    .X(_0882_));
 sky130_fd_sc_hd__inv_2 _5442_ (.A(_0882_),
    .Y(_0883_));
 sky130_fd_sc_hd__mux2_1 _5443_ (.A0(_0883_),
    .A1(_3698_),
    .S(_0870_),
    .X(_0884_));
 sky130_fd_sc_hd__inv_2 _5444_ (.A(_0884_),
    .Y(_0885_));
 sky130_fd_sc_hd__o21bai_1 _5445_ (.A1(_3589_),
    .A2(_0877_),
    .B1_N(_0000_),
    .Y(_0886_));
 sky130_fd_sc_hd__or2_1 _5446_ (.A(_0862_),
    .B(_0875_),
    .X(_0887_));
 sky130_fd_sc_hd__a22o_1 _5447_ (.A1(_0578_),
    .A2(_0885_),
    .B1(_0886_),
    .B2(_0887_),
    .X(_0888_));
 sky130_fd_sc_hd__a221o_1 _5448_ (.A1(_0855_),
    .A2(_0876_),
    .B1(_0877_),
    .B2(_0854_),
    .C1(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__o21a_1 _5449_ (.A1(_0428_),
    .A2(_1734_),
    .B1(_0571_),
    .X(_0890_));
 sky130_fd_sc_hd__nor2_1 _5450_ (.A(_0848_),
    .B(_0884_),
    .Y(_0891_));
 sky130_fd_sc_hd__o21a_1 _5451_ (.A1(_0890_),
    .A2(_0891_),
    .B1(_0575_),
    .X(_0893_));
 sky130_fd_sc_hd__a311o_1 _5452_ (.A1(_0419_),
    .A2(_0879_),
    .A3(_0880_),
    .B1(_0889_),
    .C1(_0893_),
    .X(_0894_));
 sky130_fd_sc_hd__and4b_1 _5453_ (.A_N(net140),
    .B(_0680_),
    .C(_0817_),
    .D(_0682_),
    .X(_0895_));
 sky130_fd_sc_hd__nor3_1 _5454_ (.A(_0719_),
    .B(_0810_),
    .C(_0811_),
    .Y(_0896_));
 sky130_fd_sc_hd__and2_1 _5455_ (.A(_0738_),
    .B(_0742_),
    .X(_0897_));
 sky130_fd_sc_hd__nand2_1 _5456_ (.A(_0734_),
    .B(_0735_),
    .Y(_0898_));
 sky130_fd_sc_hd__or2_1 _5457_ (.A(_0723_),
    .B(_0736_),
    .X(_0899_));
 sky130_fd_sc_hd__o211ai_2 _5458_ (.A1(_0745_),
    .A2(_0746_),
    .B1(_0764_),
    .C1(_0765_),
    .Y(_0900_));
 sky130_fd_sc_hd__a22o_1 _5459_ (.A1(_1056_),
    .A2(_0722_),
    .B1(_0875_),
    .B2(_1002_),
    .X(_0901_));
 sky130_fd_sc_hd__and4_1 _5460_ (.A(_0707_),
    .B(_0466_),
    .C(_0721_),
    .D(_0874_),
    .X(_0902_));
 sky130_fd_sc_hd__inv_2 _5461_ (.A(_0902_),
    .Y(_0904_));
 sky130_fd_sc_hd__and2_1 _5462_ (.A(_0901_),
    .B(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__or2_1 _5463_ (.A(_0727_),
    .B(_0729_),
    .X(_0906_));
 sky130_fd_sc_hd__a22oi_1 _5464_ (.A1(_0085_),
    .A2(_0325_),
    .B1(_0452_),
    .B2(_0194_),
    .Y(_0907_));
 sky130_fd_sc_hd__and4_1 _5465_ (.A(_0085_),
    .B(_1264_),
    .C(net39),
    .D(net40),
    .X(_0908_));
 sky130_fd_sc_hd__o2bb2a_1 _5466_ (.A1_N(_0739_),
    .A2_N(net41),
    .B1(_0907_),
    .B2(_0908_),
    .X(_0909_));
 sky130_fd_sc_hd__and4bb_1 _5467_ (.A_N(_0907_),
    .B_N(_0908_),
    .C(_0739_),
    .D(net41),
    .X(_0910_));
 sky130_fd_sc_hd__a211o_1 _5468_ (.A1(_0751_),
    .A2(_0752_),
    .B1(_0909_),
    .C1(_0910_),
    .X(_0911_));
 sky130_fd_sc_hd__o211ai_1 _5469_ (.A1(_0909_),
    .A2(_0910_),
    .B1(_0751_),
    .C1(_0752_),
    .Y(_0912_));
 sky130_fd_sc_hd__and2_1 _5470_ (.A(_0911_),
    .B(_0912_),
    .X(_0913_));
 sky130_fd_sc_hd__xnor2_2 _5471_ (.A(_0906_),
    .B(_0913_),
    .Y(_0915_));
 sky130_fd_sc_hd__a21bo_1 _5472_ (.A1(_0724_),
    .A2(_0732_),
    .B1_N(_0731_),
    .X(_0916_));
 sky130_fd_sc_hd__xnor2_2 _5473_ (.A(_0915_),
    .B(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__xnor2_2 _5474_ (.A(_0905_),
    .B(_0917_),
    .Y(_0918_));
 sky130_fd_sc_hd__a21oi_2 _5475_ (.A1(_0764_),
    .A2(_0900_),
    .B1(_0918_),
    .Y(_0919_));
 sky130_fd_sc_hd__and3_1 _5476_ (.A(_0764_),
    .B(_0900_),
    .C(_0918_),
    .X(_0920_));
 sky130_fd_sc_hd__a211oi_1 _5477_ (.A1(_0898_),
    .A2(_0899_),
    .B1(_0919_),
    .C1(_0920_),
    .Y(_0921_));
 sky130_fd_sc_hd__o211a_1 _5478_ (.A1(_0919_),
    .A2(_0920_),
    .B1(_0898_),
    .C1(_0899_),
    .X(_0922_));
 sky130_fd_sc_hd__and2b_1 _5479_ (.A_N(_0760_),
    .B(_0759_),
    .X(_0923_));
 sky130_fd_sc_hd__and2_2 _5480_ (.A(_0754_),
    .B(_0762_),
    .X(_0924_));
 sky130_fd_sc_hd__or3_1 _5481_ (.A(_0770_),
    .B(_0774_),
    .C(_0775_),
    .X(_0926_));
 sky130_fd_sc_hd__nand2_1 _5482_ (.A(_0769_),
    .B(_0777_),
    .Y(_0927_));
 sky130_fd_sc_hd__a22o_1 _5483_ (.A1(_2434_),
    .A2(net36),
    .B1(_0340_),
    .B2(_3442_),
    .X(_0928_));
 sky130_fd_sc_hd__nand4_4 _5484_ (.A(_3442_),
    .B(_2434_),
    .C(_0339_),
    .D(_0340_),
    .Y(_0929_));
 sky130_fd_sc_hd__nand4_2 _5485_ (.A(_2313_),
    .B(net38),
    .C(_0928_),
    .D(_0929_),
    .Y(_0930_));
 sky130_fd_sc_hd__a22o_1 _5486_ (.A1(_2324_),
    .A2(_0219_),
    .B1(_0928_),
    .B2(_0929_),
    .X(_0931_));
 sky130_fd_sc_hd__and2_1 _5487_ (.A(_0930_),
    .B(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__a22oi_1 _5488_ (.A1(_0104_),
    .A2(_3537_),
    .B1(_0105_),
    .B2(_2149_),
    .Y(_0933_));
 sky130_fd_sc_hd__and4_1 _5489_ (.A(net32),
    .B(net64),
    .C(_3537_),
    .D(_3572_),
    .X(_0934_));
 sky130_fd_sc_hd__and4bb_1 _5490_ (.A_N(_0933_),
    .B_N(_0934_),
    .C(_3644_),
    .D(_3619_),
    .X(_0935_));
 sky130_fd_sc_hd__o2bb2a_1 _5491_ (.A1_N(_3644_),
    .A2_N(_3619_),
    .B1(_0933_),
    .B2(_0934_),
    .X(_0937_));
 sky130_fd_sc_hd__nor2_1 _5492_ (.A(_0935_),
    .B(_0937_),
    .Y(_0938_));
 sky130_fd_sc_hd__o21ba_1 _5493_ (.A1(_0755_),
    .A2(_0756_),
    .B1_N(_0757_),
    .X(_0939_));
 sky130_fd_sc_hd__xnor2_2 _5494_ (.A(_0938_),
    .B(_0939_),
    .Y(_0940_));
 sky130_fd_sc_hd__xnor2_2 _5495_ (.A(_0932_),
    .B(_0940_),
    .Y(_0941_));
 sky130_fd_sc_hd__a21o_2 _5496_ (.A1(_0926_),
    .A2(_0927_),
    .B1(_0941_),
    .X(_0942_));
 sky130_fd_sc_hd__nand3_2 _5497_ (.A(_0926_),
    .B(_0927_),
    .C(_0941_),
    .Y(_0943_));
 sky130_fd_sc_hd__o211a_1 _5498_ (.A1(_0923_),
    .A2(_0924_),
    .B1(_0942_),
    .C1(_0943_),
    .X(_0944_));
 sky130_fd_sc_hd__a211oi_2 _5499_ (.A1(_0942_),
    .A2(_0943_),
    .B1(_0923_),
    .C1(_0924_),
    .Y(_0945_));
 sky130_fd_sc_hd__nand3_2 _5500_ (.A(_0778_),
    .B(_0797_),
    .C(_0798_),
    .Y(_0946_));
 sky130_fd_sc_hd__or2_1 _5501_ (.A(_0773_),
    .B(_0774_),
    .X(_0948_));
 sky130_fd_sc_hd__a32o_1 _5502_ (.A1(_2892_),
    .A2(_2707_),
    .A3(_0781_),
    .B1(_0780_),
    .B2(_2773_),
    .X(_0949_));
 sky130_fd_sc_hd__a22o_1 _5503_ (.A1(_3431_),
    .A2(net4),
    .B1(net5),
    .B2(_3433_),
    .X(_0950_));
 sky130_fd_sc_hd__nand4_1 _5504_ (.A(_3195_),
    .B(_3633_),
    .C(_2642_),
    .D(_2686_),
    .Y(_0951_));
 sky130_fd_sc_hd__a22oi_1 _5505_ (.A1(_3631_),
    .A2(_2248_),
    .B1(_0950_),
    .B2(_0951_),
    .Y(_0952_));
 sky130_fd_sc_hd__and4_1 _5506_ (.A(_3343_),
    .B(_2248_),
    .C(_0950_),
    .D(_0951_),
    .X(_0953_));
 sky130_fd_sc_hd__or2_1 _5507_ (.A(_0952_),
    .B(_0953_),
    .X(_0954_));
 sky130_fd_sc_hd__xnor2_1 _5508_ (.A(_0949_),
    .B(_0954_),
    .Y(_0955_));
 sky130_fd_sc_hd__xor2_1 _5509_ (.A(_0948_),
    .B(_0955_),
    .X(_0956_));
 sky130_fd_sc_hd__nand2_1 _5510_ (.A(_2881_),
    .B(_2751_),
    .Y(_0957_));
 sky130_fd_sc_hd__and3_1 _5511_ (.A(_3352_),
    .B(_0373_),
    .C(net7),
    .X(_0959_));
 sky130_fd_sc_hd__a22o_1 _5512_ (.A1(_0373_),
    .A2(net7),
    .B1(net8),
    .B2(_3352_),
    .X(_0960_));
 sky130_fd_sc_hd__a21bo_1 _5513_ (.A1(_2489_),
    .A2(_0959_),
    .B1_N(_0960_),
    .X(_0961_));
 sky130_fd_sc_hd__xor2_2 _5514_ (.A(_0957_),
    .B(_0961_),
    .X(_0962_));
 sky130_fd_sc_hd__and2_1 _5515_ (.A(_0281_),
    .B(_2521_),
    .X(_0963_));
 sky130_fd_sc_hd__a22o_1 _5516_ (.A1(_0390_),
    .A2(net10),
    .B1(net11),
    .B2(_0488_),
    .X(_0964_));
 sky130_fd_sc_hd__nand4_2 _5517_ (.A(_3451_),
    .B(_3448_),
    .C(_2565_),
    .D(_2598_),
    .Y(_0965_));
 sky130_fd_sc_hd__nand3_1 _5518_ (.A(_0963_),
    .B(_0964_),
    .C(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__a21o_1 _5519_ (.A1(_0964_),
    .A2(_0965_),
    .B1(_0963_),
    .X(_0967_));
 sky130_fd_sc_hd__a21bo_1 _5520_ (.A1(_0785_),
    .A2(_0786_),
    .B1_N(_0787_),
    .X(_0968_));
 sky130_fd_sc_hd__nand3_1 _5521_ (.A(_0966_),
    .B(_0967_),
    .C(_0968_),
    .Y(_0970_));
 sky130_fd_sc_hd__a21o_1 _5522_ (.A1(_0966_),
    .A2(_0967_),
    .B1(_0968_),
    .X(_0971_));
 sky130_fd_sc_hd__nand3_2 _5523_ (.A(_0962_),
    .B(_0970_),
    .C(_0971_),
    .Y(_0972_));
 sky130_fd_sc_hd__a21o_1 _5524_ (.A1(_0970_),
    .A2(_0971_),
    .B1(_0962_),
    .X(_0973_));
 sky130_fd_sc_hd__a21bo_1 _5525_ (.A1(_0784_),
    .A2(_0792_),
    .B1_N(_0791_),
    .X(_0974_));
 sky130_fd_sc_hd__nand3_4 _5526_ (.A(_0972_),
    .B(_0973_),
    .C(_0974_),
    .Y(_0975_));
 sky130_fd_sc_hd__a21o_1 _5527_ (.A1(_0972_),
    .A2(_0973_),
    .B1(_0974_),
    .X(_0976_));
 sky130_fd_sc_hd__and3_1 _5528_ (.A(_0956_),
    .B(_0975_),
    .C(_0976_),
    .X(_0977_));
 sky130_fd_sc_hd__a21oi_2 _5529_ (.A1(_0975_),
    .A2(_0976_),
    .B1(_0956_),
    .Y(_0978_));
 sky130_fd_sc_hd__a211oi_4 _5530_ (.A1(_0797_),
    .A2(_0946_),
    .B1(_0977_),
    .C1(_0978_),
    .Y(_0979_));
 sky130_fd_sc_hd__o211a_1 _5531_ (.A1(_0977_),
    .A2(_0978_),
    .B1(_0797_),
    .C1(_0946_),
    .X(_0981_));
 sky130_fd_sc_hd__or4_2 _5532_ (.A(_0944_),
    .B(_0945_),
    .C(_0979_),
    .D(_0981_),
    .X(_0982_));
 sky130_fd_sc_hd__o22ai_2 _5533_ (.A1(_0944_),
    .A2(_0945_),
    .B1(_0979_),
    .B2(_0981_),
    .Y(_0983_));
 sky130_fd_sc_hd__o211a_1 _5534_ (.A1(_0801_),
    .A2(_0803_),
    .B1(_0982_),
    .C1(_0983_),
    .X(_0984_));
 sky130_fd_sc_hd__a211oi_2 _5535_ (.A1(_0982_),
    .A2(_0983_),
    .B1(_0801_),
    .C1(_0803_),
    .Y(_0985_));
 sky130_fd_sc_hd__nor4_1 _5536_ (.A(_0921_),
    .B(_0922_),
    .C(_0984_),
    .D(_0985_),
    .Y(_0986_));
 sky130_fd_sc_hd__o22a_1 _5537_ (.A1(_0921_),
    .A2(_0922_),
    .B1(_0984_),
    .B2(_0985_),
    .X(_0987_));
 sky130_fd_sc_hd__a211oi_1 _5538_ (.A1(_0806_),
    .A2(_0808_),
    .B1(net106),
    .C1(_0987_),
    .Y(_0988_));
 sky130_fd_sc_hd__o211a_1 _5539_ (.A1(net106),
    .A2(_0987_),
    .B1(_0806_),
    .C1(_0808_),
    .X(_0989_));
 sky130_fd_sc_hd__or3_1 _5540_ (.A(_0897_),
    .B(_0988_),
    .C(_0989_),
    .X(_0990_));
 sky130_fd_sc_hd__o21ai_1 _5541_ (.A1(_0988_),
    .A2(_0989_),
    .B1(_0897_),
    .Y(_0992_));
 sky130_fd_sc_hd__o211a_1 _5542_ (.A1(_0810_),
    .A2(_0896_),
    .B1(_0990_),
    .C1(_0992_),
    .X(_0993_));
 sky130_fd_sc_hd__a211o_1 _5543_ (.A1(_0990_),
    .A2(_0992_),
    .B1(_0810_),
    .C1(_0896_),
    .X(_0994_));
 sky130_fd_sc_hd__or2b_1 _5544_ (.A(_0993_),
    .B_N(_0994_),
    .X(_0995_));
 sky130_fd_sc_hd__a21o_1 _5545_ (.A1(net140),
    .A2(_0815_),
    .B1(_0814_),
    .X(_0996_));
 sky130_fd_sc_hd__xnor2_1 _5546_ (.A(_0995_),
    .B(_0996_),
    .Y(_0997_));
 sky130_fd_sc_hd__o21ai_1 _5547_ (.A1(_0824_),
    .A2(_0895_),
    .B1(_0997_),
    .Y(_0998_));
 sky130_fd_sc_hd__or3_1 _5548_ (.A(_0824_),
    .B(_0997_),
    .C(_0895_),
    .X(_0999_));
 sky130_fd_sc_hd__and2b_1 _5549_ (.A_N(_0722_),
    .B(_2587_),
    .X(_1000_));
 sky130_fd_sc_hd__a21o_1 _5550_ (.A1(_0829_),
    .A2(_0831_),
    .B1(_1000_),
    .X(_1001_));
 sky130_fd_sc_hd__a21oi_1 _5551_ (.A1(_0878_),
    .A2(_1001_),
    .B1(_0181_),
    .Y(_1003_));
 sky130_fd_sc_hd__o21a_1 _5552_ (.A1(_0878_),
    .A2(_1001_),
    .B1(_1003_),
    .X(_1004_));
 sky130_fd_sc_hd__a31o_1 _5553_ (.A1(_0320_),
    .A2(_0998_),
    .A3(_0999_),
    .B1(_1004_),
    .X(_1005_));
 sky130_fd_sc_hd__or3_1 _5554_ (.A(_0872_),
    .B(_0894_),
    .C(_1005_),
    .X(_1006_));
 sky130_fd_sc_hd__clkbuf_4 _5555_ (.A(_1006_),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_4 _5556_ (.A(net45),
    .X(_1007_));
 sky130_fd_sc_hd__clkbuf_4 _5557_ (.A(_1007_),
    .X(_1008_));
 sky130_fd_sc_hd__nor2_1 _5558_ (.A(_1876_),
    .B(_1008_),
    .Y(_1009_));
 sky130_fd_sc_hd__and2_1 _5559_ (.A(_1876_),
    .B(_1008_),
    .X(_1010_));
 sky130_fd_sc_hd__or2_2 _5560_ (.A(_1009_),
    .B(_1010_),
    .X(_1011_));
 sky130_fd_sc_hd__and2b_1 _5561_ (.A_N(_0875_),
    .B(_0862_),
    .X(_1013_));
 sky130_fd_sc_hd__a21o_1 _5562_ (.A1(_0878_),
    .A2(_1001_),
    .B1(_1013_),
    .X(_1014_));
 sky130_fd_sc_hd__or2_1 _5563_ (.A(_1011_),
    .B(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__a21oi_1 _5564_ (.A1(_1011_),
    .A2(_1014_),
    .B1(_0181_),
    .Y(_1016_));
 sky130_fd_sc_hd__mux4_1 _5565_ (.A0(_1876_),
    .A1(_0862_),
    .A2(_2587_),
    .A3(_3128_),
    .S0(_0583_),
    .S1(_0584_),
    .X(_1017_));
 sky130_fd_sc_hd__mux2_1 _5566_ (.A0(_0585_),
    .A1(_1017_),
    .S(_0429_),
    .X(_1018_));
 sky130_fd_sc_hd__o2bb2a_1 _5567_ (.A1_N(_0428_),
    .A2_N(_1122_),
    .B1(_0005_),
    .B2(_0189_),
    .X(_1019_));
 sky130_fd_sc_hd__o311a_1 _5568_ (.A1(_0199_),
    .A2(_0848_),
    .A3(_1018_),
    .B1(_1019_),
    .C1(_0849_),
    .X(_1020_));
 sky130_fd_sc_hd__nand2_1 _5569_ (.A(_1876_),
    .B(_1008_),
    .Y(_1021_));
 sky130_fd_sc_hd__a21oi_1 _5570_ (.A1(_0438_),
    .A2(_1021_),
    .B1(_0000_),
    .Y(_1022_));
 sky130_fd_sc_hd__nor2_1 _5571_ (.A(_1009_),
    .B(_1022_),
    .Y(_1024_));
 sky130_fd_sc_hd__a221o_1 _5572_ (.A1(_0855_),
    .A2(_1009_),
    .B1(_1010_),
    .B2(_0854_),
    .C1(_1024_),
    .X(_1025_));
 sky130_fd_sc_hd__a211o_1 _5573_ (.A1(_2095_),
    .A2(_0578_),
    .B1(_1020_),
    .C1(_1025_),
    .X(_1026_));
 sky130_fd_sc_hd__o31ai_4 _5574_ (.A1(_0826_),
    .A2(_0836_),
    .A3(_0877_),
    .B1(_0887_),
    .Y(_1027_));
 sky130_fd_sc_hd__nand2_1 _5575_ (.A(_1011_),
    .B(_1027_),
    .Y(_1028_));
 sky130_fd_sc_hd__or2_1 _5576_ (.A(_1011_),
    .B(_1027_),
    .X(_1029_));
 sky130_fd_sc_hd__a21o_1 _5577_ (.A1(_0573_),
    .A2(_2095_),
    .B1(_0890_),
    .X(_1030_));
 sky130_fd_sc_hd__a32o_1 _5578_ (.A1(_0419_),
    .A2(_1028_),
    .A3(_1029_),
    .B1(_1030_),
    .B2(_0575_),
    .X(_1031_));
 sky130_fd_sc_hd__or2_1 _5579_ (.A(_1026_),
    .B(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__inv_2 _5580_ (.A(_0919_),
    .Y(_1033_));
 sky130_fd_sc_hd__a211o_1 _5581_ (.A1(_0898_),
    .A2(_0899_),
    .B1(_0919_),
    .C1(_0920_),
    .X(_1035_));
 sky130_fd_sc_hd__and2b_1 _5582_ (.A_N(_0915_),
    .B(_0916_),
    .X(_1036_));
 sky130_fd_sc_hd__a21oi_1 _5583_ (.A1(_0905_),
    .A2(_0917_),
    .B1(_1036_),
    .Y(_1037_));
 sky130_fd_sc_hd__o211ai_4 _5584_ (.A1(_0923_),
    .A2(_0924_),
    .B1(_0942_),
    .C1(_0943_),
    .Y(_1038_));
 sky130_fd_sc_hd__a22o_1 _5585_ (.A1(_0335_),
    .A2(_0720_),
    .B1(_0873_),
    .B2(_0434_),
    .X(_1039_));
 sky130_fd_sc_hd__nand4_1 _5586_ (.A(_0335_),
    .B(_0434_),
    .C(_0721_),
    .D(_0874_),
    .Y(_1040_));
 sky130_fd_sc_hd__nand2_1 _5587_ (.A(_1039_),
    .B(_1040_),
    .Y(_1041_));
 sky130_fd_sc_hd__nand2_1 _5588_ (.A(_0466_),
    .B(_1007_),
    .Y(_1042_));
 sky130_fd_sc_hd__xnor2_1 _5589_ (.A(_1041_),
    .B(_1042_),
    .Y(_1043_));
 sky130_fd_sc_hd__nor2_1 _5590_ (.A(_0904_),
    .B(_1043_),
    .Y(_1044_));
 sky130_fd_sc_hd__and2_1 _5591_ (.A(_0904_),
    .B(_1043_),
    .X(_1046_));
 sky130_fd_sc_hd__or2_1 _5592_ (.A(_1044_),
    .B(_1046_),
    .X(_1047_));
 sky130_fd_sc_hd__nand2_1 _5593_ (.A(_0906_),
    .B(_0913_),
    .Y(_1048_));
 sky130_fd_sc_hd__or2_1 _5594_ (.A(_0908_),
    .B(_0910_),
    .X(_1049_));
 sky130_fd_sc_hd__a22oi_1 _5595_ (.A1(_3635_),
    .A2(_0325_),
    .B1(_0452_),
    .B2(_3440_),
    .Y(_1050_));
 sky130_fd_sc_hd__and4_1 _5596_ (.A(_0085_),
    .B(_2302_),
    .C(_0325_),
    .D(_0452_),
    .X(_1051_));
 sky130_fd_sc_hd__o2bb2a_1 _5597_ (.A1_N(_1275_),
    .A2_N(_0654_),
    .B1(_1050_),
    .B2(_1051_),
    .X(_1052_));
 sky130_fd_sc_hd__and4bb_1 _5598_ (.A_N(_1050_),
    .B_N(_1051_),
    .C(_1275_),
    .D(net41),
    .X(_1053_));
 sky130_fd_sc_hd__a211o_1 _5599_ (.A1(_0929_),
    .A2(_0930_),
    .B1(_1052_),
    .C1(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__o211ai_1 _5600_ (.A1(_1052_),
    .A2(_1053_),
    .B1(_0929_),
    .C1(_0930_),
    .Y(_1055_));
 sky130_fd_sc_hd__and2_1 _5601_ (.A(_1054_),
    .B(_1055_),
    .X(_1057_));
 sky130_fd_sc_hd__xnor2_1 _5602_ (.A(_1049_),
    .B(_1057_),
    .Y(_1058_));
 sky130_fd_sc_hd__a21oi_1 _5603_ (.A1(_0911_),
    .A2(_1048_),
    .B1(_1058_),
    .Y(_1059_));
 sky130_fd_sc_hd__and3_1 _5604_ (.A(_0911_),
    .B(_1048_),
    .C(_1058_),
    .X(_1060_));
 sky130_fd_sc_hd__nor3_1 _5605_ (.A(_1047_),
    .B(_1059_),
    .C(_1060_),
    .Y(_1061_));
 sky130_fd_sc_hd__o21a_1 _5606_ (.A1(_1059_),
    .A2(_1060_),
    .B1(_1047_),
    .X(_1062_));
 sky130_fd_sc_hd__a211oi_2 _5607_ (.A1(_0942_),
    .A2(_1038_),
    .B1(_1061_),
    .C1(_1062_),
    .Y(_1063_));
 sky130_fd_sc_hd__o211a_1 _5608_ (.A1(_1061_),
    .A2(_1062_),
    .B1(_0942_),
    .C1(_1038_),
    .X(_1064_));
 sky130_fd_sc_hd__nor3_2 _5609_ (.A(_1037_),
    .B(_1063_),
    .C(_1064_),
    .Y(_1065_));
 sky130_fd_sc_hd__o21a_1 _5610_ (.A1(_1063_),
    .A2(_1064_),
    .B1(_1037_),
    .X(_1066_));
 sky130_fd_sc_hd__nor4_1 _5611_ (.A(_0944_),
    .B(_0945_),
    .C(_0979_),
    .D(_0981_),
    .Y(_1068_));
 sky130_fd_sc_hd__nand2_1 _5612_ (.A(_0932_),
    .B(_0940_),
    .Y(_1069_));
 sky130_fd_sc_hd__o31a_1 _5613_ (.A1(_0935_),
    .A2(_0937_),
    .A3(_0939_),
    .B1(_1069_),
    .X(_1070_));
 sky130_fd_sc_hd__and2b_1 _5614_ (.A_N(_0954_),
    .B(_0949_),
    .X(_1071_));
 sky130_fd_sc_hd__and2_1 _5615_ (.A(_0948_),
    .B(_0955_),
    .X(_1072_));
 sky130_fd_sc_hd__a22o_1 _5616_ (.A1(_3644_),
    .A2(_0339_),
    .B1(_0340_),
    .B2(_2434_),
    .X(_1073_));
 sky130_fd_sc_hd__nand4_4 _5617_ (.A(_2434_),
    .B(_3644_),
    .C(_0339_),
    .D(_0340_),
    .Y(_1074_));
 sky130_fd_sc_hd__a22o_1 _5618_ (.A1(_2390_),
    .A2(_0220_),
    .B1(_1073_),
    .B2(_1074_),
    .X(_1075_));
 sky130_fd_sc_hd__nand4_2 _5619_ (.A(_2390_),
    .B(_0219_),
    .C(_1073_),
    .D(_1074_),
    .Y(_1076_));
 sky130_fd_sc_hd__nand2_1 _5620_ (.A(_1075_),
    .B(_1076_),
    .Y(_1077_));
 sky130_fd_sc_hd__nand2_1 _5621_ (.A(_3422_),
    .B(_3651_),
    .Y(_1079_));
 sky130_fd_sc_hd__xnor2_1 _5622_ (.A(_3573_),
    .B(_1079_),
    .Y(_1080_));
 sky130_fd_sc_hd__nand2_1 _5623_ (.A(_2160_),
    .B(_0110_),
    .Y(_1081_));
 sky130_fd_sc_hd__xnor2_1 _5624_ (.A(_1080_),
    .B(_1081_),
    .Y(_1082_));
 sky130_fd_sc_hd__nor2_1 _5625_ (.A(_0934_),
    .B(_0935_),
    .Y(_1083_));
 sky130_fd_sc_hd__xor2_1 _5626_ (.A(_1082_),
    .B(_1083_),
    .X(_1084_));
 sky130_fd_sc_hd__xor2_1 _5627_ (.A(_1077_),
    .B(_1084_),
    .X(_1085_));
 sky130_fd_sc_hd__o21a_1 _5628_ (.A1(_1071_),
    .A2(_1072_),
    .B1(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__nor3_1 _5629_ (.A(_1071_),
    .B(_1072_),
    .C(_1085_),
    .Y(_1087_));
 sky130_fd_sc_hd__nor3_1 _5630_ (.A(_1070_),
    .B(_1086_),
    .C(_1087_),
    .Y(_1088_));
 sky130_fd_sc_hd__o21a_1 _5631_ (.A1(_1086_),
    .A2(_1087_),
    .B1(_1070_),
    .X(_1090_));
 sky130_fd_sc_hd__nand3_1 _5632_ (.A(_0956_),
    .B(_0975_),
    .C(_0976_),
    .Y(_1091_));
 sky130_fd_sc_hd__a41o_1 _5633_ (.A1(_3197_),
    .A2(_3272_),
    .A3(_2664_),
    .A4(_2707_),
    .B1(_0953_),
    .X(_1092_));
 sky130_fd_sc_hd__a32o_1 _5634_ (.A1(_2892_),
    .A2(_2751_),
    .A3(_0960_),
    .B1(_0959_),
    .B2(_2499_),
    .X(_1093_));
 sky130_fd_sc_hd__a22o_1 _5635_ (.A1(net162),
    .A2(net5),
    .B1(net6),
    .B2(_3433_),
    .X(_1094_));
 sky130_fd_sc_hd__nand4_1 _5636_ (.A(_3195_),
    .B(_3431_),
    .C(net5),
    .D(net6),
    .Y(_1095_));
 sky130_fd_sc_hd__a22oi_1 _5637_ (.A1(_3430_),
    .A2(_0491_),
    .B1(_1094_),
    .B2(_1095_),
    .Y(_1096_));
 sky130_fd_sc_hd__and4_1 _5638_ (.A(_3343_),
    .B(_0491_),
    .C(_1094_),
    .D(_1095_),
    .X(_1097_));
 sky130_fd_sc_hd__or2_1 _5639_ (.A(_1096_),
    .B(_1097_),
    .X(_1098_));
 sky130_fd_sc_hd__xnor2_1 _5640_ (.A(_1093_),
    .B(_1098_),
    .Y(_1099_));
 sky130_fd_sc_hd__xnor2_1 _5641_ (.A(_1092_),
    .B(_1099_),
    .Y(_1101_));
 sky130_fd_sc_hd__and3_1 _5642_ (.A(_3352_),
    .B(_0373_),
    .C(net8),
    .X(_1102_));
 sky130_fd_sc_hd__a22o_1 _5643_ (.A1(_0373_),
    .A2(net8),
    .B1(net9),
    .B2(_3352_),
    .X(_1103_));
 sky130_fd_sc_hd__a21bo_1 _5644_ (.A1(_2532_),
    .A2(_1102_),
    .B1_N(_1103_),
    .X(_1104_));
 sky130_fd_sc_hd__nand2_1 _5645_ (.A(_0042_),
    .B(_2773_),
    .Y(_1105_));
 sky130_fd_sc_hd__xor2_1 _5646_ (.A(_1104_),
    .B(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__and2_1 _5647_ (.A(_0281_),
    .B(net10),
    .X(_1107_));
 sky130_fd_sc_hd__nand4_1 _5648_ (.A(_3451_),
    .B(_3452_),
    .C(_2598_),
    .D(_1854_),
    .Y(_1108_));
 sky130_fd_sc_hd__a22o_1 _5649_ (.A1(_0390_),
    .A2(net11),
    .B1(_1854_),
    .B2(_0488_),
    .X(_1109_));
 sky130_fd_sc_hd__nand3_1 _5650_ (.A(_1107_),
    .B(_1108_),
    .C(_1109_),
    .Y(_1110_));
 sky130_fd_sc_hd__a21o_1 _5651_ (.A1(_1108_),
    .A2(_1109_),
    .B1(_1107_),
    .X(_1112_));
 sky130_fd_sc_hd__a21bo_1 _5652_ (.A1(_0963_),
    .A2(_0964_),
    .B1_N(_0965_),
    .X(_1113_));
 sky130_fd_sc_hd__nand3_1 _5653_ (.A(_1110_),
    .B(_1112_),
    .C(_1113_),
    .Y(_1114_));
 sky130_fd_sc_hd__a21o_1 _5654_ (.A1(_1110_),
    .A2(_1112_),
    .B1(_1113_),
    .X(_1115_));
 sky130_fd_sc_hd__nand3_1 _5655_ (.A(_1106_),
    .B(_1114_),
    .C(_1115_),
    .Y(_1116_));
 sky130_fd_sc_hd__a21o_1 _5656_ (.A1(_1114_),
    .A2(_1115_),
    .B1(_1106_),
    .X(_1117_));
 sky130_fd_sc_hd__a21bo_1 _5657_ (.A1(_0962_),
    .A2(_0971_),
    .B1_N(_0970_),
    .X(_1118_));
 sky130_fd_sc_hd__and3_2 _5658_ (.A(_1116_),
    .B(_1117_),
    .C(_1118_),
    .X(_1119_));
 sky130_fd_sc_hd__a21oi_2 _5659_ (.A1(_1116_),
    .A2(_1117_),
    .B1(_1118_),
    .Y(_1120_));
 sky130_fd_sc_hd__nor3_2 _5660_ (.A(_1101_),
    .B(_1119_),
    .C(_1120_),
    .Y(_1121_));
 sky130_fd_sc_hd__o21a_1 _5661_ (.A1(_1119_),
    .A2(_1120_),
    .B1(_1101_),
    .X(_1123_));
 sky130_fd_sc_hd__a211o_2 _5662_ (.A1(_0975_),
    .A2(_1091_),
    .B1(_1121_),
    .C1(_1123_),
    .X(_1124_));
 sky130_fd_sc_hd__o211ai_2 _5663_ (.A1(_1121_),
    .A2(_1123_),
    .B1(_0975_),
    .C1(_1091_),
    .Y(_1125_));
 sky130_fd_sc_hd__or4bb_2 _5664_ (.A(net118),
    .B(_1090_),
    .C_N(_1124_),
    .D_N(_1125_),
    .X(_1126_));
 sky130_fd_sc_hd__a2bb2o_1 _5665_ (.A1_N(_1088_),
    .A2_N(_1090_),
    .B1(_1124_),
    .B2(_1125_),
    .X(_1127_));
 sky130_fd_sc_hd__o211a_2 _5666_ (.A1(net119),
    .A2(net111),
    .B1(_1126_),
    .C1(_1127_),
    .X(_1128_));
 sky130_fd_sc_hd__a211oi_4 _5667_ (.A1(net136),
    .A2(_1127_),
    .B1(net119),
    .C1(net110),
    .Y(_1129_));
 sky130_fd_sc_hd__or4_2 _5668_ (.A(_1065_),
    .B(_1066_),
    .C(_1128_),
    .D(_1129_),
    .X(_1130_));
 sky130_fd_sc_hd__o22ai_4 _5669_ (.A1(_1065_),
    .A2(_1066_),
    .B1(_1128_),
    .B2(_1129_),
    .Y(_1131_));
 sky130_fd_sc_hd__o211a_1 _5670_ (.A1(net130),
    .A2(net106),
    .B1(_1130_),
    .C1(_1131_),
    .X(_1132_));
 sky130_fd_sc_hd__a211oi_1 _5671_ (.A1(_1130_),
    .A2(_1131_),
    .B1(net130),
    .C1(net106),
    .Y(_1134_));
 sky130_fd_sc_hd__a211o_1 _5672_ (.A1(_1033_),
    .A2(_1035_),
    .B1(_1132_),
    .C1(_1134_),
    .X(_1135_));
 sky130_fd_sc_hd__o211ai_2 _5673_ (.A1(_1132_),
    .A2(net161),
    .B1(_1033_),
    .C1(_1035_),
    .Y(_1136_));
 sky130_fd_sc_hd__o21bai_1 _5674_ (.A1(_0897_),
    .A2(_0989_),
    .B1_N(_0988_),
    .Y(_1137_));
 sky130_fd_sc_hd__nand3_2 _5675_ (.A(net134),
    .B(_1136_),
    .C(_1137_),
    .Y(_1138_));
 sky130_fd_sc_hd__a21o_1 _5676_ (.A1(_1135_),
    .A2(_1136_),
    .B1(_1137_),
    .X(_1139_));
 sky130_fd_sc_hd__nand2_1 _5677_ (.A(_1138_),
    .B(_1139_),
    .Y(_1140_));
 sky130_fd_sc_hd__a21oi_1 _5678_ (.A1(_0814_),
    .A2(_0994_),
    .B1(_0993_),
    .Y(_1141_));
 sky130_fd_sc_hd__xnor2_1 _5679_ (.A(_1140_),
    .B(_1141_),
    .Y(_1142_));
 sky130_fd_sc_hd__or2b_1 _5680_ (.A(_0819_),
    .B_N(_0997_),
    .X(_1143_));
 sky130_fd_sc_hd__or2_1 _5681_ (.A(_0821_),
    .B(_1143_),
    .X(_1145_));
 sky130_fd_sc_hd__a31o_1 _5682_ (.A1(_0549_),
    .A2(net164),
    .A3(_0553_),
    .B1(_1145_),
    .X(_1146_));
 sky130_fd_sc_hd__nand2_1 _5683_ (.A(net141),
    .B(_0817_),
    .Y(_1147_));
 sky130_fd_sc_hd__nand2_1 _5684_ (.A(_0997_),
    .B(_0895_),
    .Y(_1148_));
 sky130_fd_sc_hd__o221a_1 _5685_ (.A1(_0995_),
    .A2(_1147_),
    .B1(_1143_),
    .B2(_0820_),
    .C1(_1148_),
    .X(_1149_));
 sky130_fd_sc_hd__nand3_1 _5686_ (.A(_1142_),
    .B(_1146_),
    .C(_1149_),
    .Y(_1150_));
 sky130_fd_sc_hd__a21o_1 _5687_ (.A1(_1146_),
    .A2(_1149_),
    .B1(_1142_),
    .X(_1151_));
 sky130_fd_sc_hd__and3_1 _5688_ (.A(_0320_),
    .B(_1150_),
    .C(_1151_),
    .X(_1152_));
 sky130_fd_sc_hd__a211o_2 _5689_ (.A1(_1015_),
    .A2(_1016_),
    .B1(_1032_),
    .C1(_1152_),
    .X(net81));
 sky130_fd_sc_hd__inv_2 _5690_ (.A(_0814_),
    .Y(_1153_));
 sky130_fd_sc_hd__or3_2 _5691_ (.A(_1153_),
    .B(_0995_),
    .C(_1140_),
    .X(_1155_));
 sky130_fd_sc_hd__nor2_1 _5692_ (.A(_1063_),
    .B(_1065_),
    .Y(_1156_));
 sky130_fd_sc_hd__xnor2_1 _5693_ (.A(_1044_),
    .B(_1156_),
    .Y(_1157_));
 sky130_fd_sc_hd__nor4_1 _5694_ (.A(_1065_),
    .B(_1066_),
    .C(_1128_),
    .D(_1129_),
    .Y(_1158_));
 sky130_fd_sc_hd__nor2_1 _5695_ (.A(_1059_),
    .B(_1061_),
    .Y(_1159_));
 sky130_fd_sc_hd__and4_1 _5696_ (.A(_1264_),
    .B(_0314_),
    .C(net42),
    .D(net43),
    .X(_1160_));
 sky130_fd_sc_hd__inv_2 _5697_ (.A(_1160_),
    .Y(_1161_));
 sky130_fd_sc_hd__a22o_1 _5698_ (.A1(_1275_),
    .A2(_0720_),
    .B1(_0873_),
    .B2(_0739_),
    .X(_1162_));
 sky130_fd_sc_hd__and4_1 _5699_ (.A(_0434_),
    .B(net45),
    .C(_1161_),
    .D(_1162_),
    .X(_1163_));
 sky130_fd_sc_hd__a22oi_1 _5700_ (.A1(_0707_),
    .A2(_1007_),
    .B1(_1161_),
    .B2(_1162_),
    .Y(_1164_));
 sky130_fd_sc_hd__or2_1 _5701_ (.A(_1163_),
    .B(_1164_),
    .X(_1166_));
 sky130_fd_sc_hd__o21ai_2 _5702_ (.A1(_1041_),
    .A2(_1042_),
    .B1(_1040_),
    .Y(_1167_));
 sky130_fd_sc_hd__xnor2_2 _5703_ (.A(_1166_),
    .B(_1167_),
    .Y(_1168_));
 sky130_fd_sc_hd__clkbuf_4 _5704_ (.A(net46),
    .X(_1169_));
 sky130_fd_sc_hd__buf_4 _5705_ (.A(_1169_),
    .X(_1170_));
 sky130_fd_sc_hd__nand2_1 _5706_ (.A(_1002_),
    .B(_1170_),
    .Y(_1171_));
 sky130_fd_sc_hd__xnor2_2 _5707_ (.A(_1168_),
    .B(_1171_),
    .Y(_1172_));
 sky130_fd_sc_hd__nand2_1 _5708_ (.A(_1049_),
    .B(_1057_),
    .Y(_1173_));
 sky130_fd_sc_hd__or2_1 _5709_ (.A(_1051_),
    .B(_1053_),
    .X(_1174_));
 sky130_fd_sc_hd__and4_1 _5710_ (.A(_3635_),
    .B(_3442_),
    .C(_0325_),
    .D(_0452_),
    .X(_1175_));
 sky130_fd_sc_hd__a22oi_1 _5711_ (.A1(_3442_),
    .A2(_0326_),
    .B1(_0453_),
    .B2(_3635_),
    .Y(_1177_));
 sky130_fd_sc_hd__and4bb_1 _5712_ (.A_N(_1175_),
    .B_N(_1177_),
    .C(_0095_),
    .D(_0654_),
    .X(_1178_));
 sky130_fd_sc_hd__o2bb2a_1 _5713_ (.A1_N(_0095_),
    .A2_N(_0654_),
    .B1(_1175_),
    .B2(_1177_),
    .X(_1179_));
 sky130_fd_sc_hd__a211o_1 _5714_ (.A1(_1074_),
    .A2(_1076_),
    .B1(_1178_),
    .C1(_1179_),
    .X(_1180_));
 sky130_fd_sc_hd__o211ai_1 _5715_ (.A1(_1178_),
    .A2(_1179_),
    .B1(_1074_),
    .C1(_1076_),
    .Y(_1181_));
 sky130_fd_sc_hd__and2_1 _5716_ (.A(_1180_),
    .B(_1181_),
    .X(_1182_));
 sky130_fd_sc_hd__xnor2_1 _5717_ (.A(_1174_),
    .B(_1182_),
    .Y(_1183_));
 sky130_fd_sc_hd__a21o_1 _5718_ (.A1(_1054_),
    .A2(_1173_),
    .B1(_1183_),
    .X(_1184_));
 sky130_fd_sc_hd__nand3_1 _5719_ (.A(_1054_),
    .B(_1173_),
    .C(_1183_),
    .Y(_1185_));
 sky130_fd_sc_hd__nand3_2 _5720_ (.A(_1172_),
    .B(_1184_),
    .C(_1185_),
    .Y(_1186_));
 sky130_fd_sc_hd__a21o_1 _5721_ (.A1(_1184_),
    .A2(_1185_),
    .B1(_1172_),
    .X(_1188_));
 sky130_fd_sc_hd__o211a_1 _5722_ (.A1(net187),
    .A2(net118),
    .B1(_1186_),
    .C1(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__a211oi_1 _5723_ (.A1(_1186_),
    .A2(_1188_),
    .B1(net187),
    .C1(net118),
    .Y(_1190_));
 sky130_fd_sc_hd__nor3_1 _5724_ (.A(_1159_),
    .B(_1189_),
    .C(_1190_),
    .Y(_1191_));
 sky130_fd_sc_hd__o21a_1 _5725_ (.A1(_1189_),
    .A2(_1190_),
    .B1(_1159_),
    .X(_1192_));
 sky130_fd_sc_hd__or2b_1 _5726_ (.A(_1083_),
    .B_N(_1082_),
    .X(_1193_));
 sky130_fd_sc_hd__or2_2 _5727_ (.A(_1077_),
    .B(_1084_),
    .X(_1194_));
 sky130_fd_sc_hd__and2b_1 _5728_ (.A_N(_1098_),
    .B(_1093_),
    .X(_1195_));
 sky130_fd_sc_hd__and2_1 _5729_ (.A(_1092_),
    .B(_1099_),
    .X(_1196_));
 sky130_fd_sc_hd__nand4_4 _5730_ (.A(_2106_),
    .B(_2149_),
    .C(_0339_),
    .D(_0340_),
    .Y(_1197_));
 sky130_fd_sc_hd__a22o_1 _5731_ (.A1(_2149_),
    .A2(net36),
    .B1(net37),
    .B2(_2106_),
    .X(_1199_));
 sky130_fd_sc_hd__nand4_2 _5732_ (.A(_3530_),
    .B(net38),
    .C(_1197_),
    .D(_1199_),
    .Y(_1200_));
 sky130_fd_sc_hd__a22o_1 _5733_ (.A1(_2445_),
    .A2(_0220_),
    .B1(_1197_),
    .B2(_1199_),
    .X(_1201_));
 sky130_fd_sc_hd__nand2_1 _5734_ (.A(_1200_),
    .B(_1201_),
    .Y(_1202_));
 sky130_fd_sc_hd__and4_1 _5735_ (.A(net64),
    .B(_3572_),
    .C(net3),
    .D(_2642_),
    .X(_1203_));
 sky130_fd_sc_hd__a22o_1 _5736_ (.A1(_3572_),
    .A2(_3651_),
    .B1(_2642_),
    .B2(_3422_),
    .X(_1204_));
 sky130_fd_sc_hd__or2b_1 _5737_ (.A(_1203_),
    .B_N(_1204_),
    .X(_1205_));
 sky130_fd_sc_hd__nand2_1 _5738_ (.A(_2215_),
    .B(_0110_),
    .Y(_1206_));
 sky130_fd_sc_hd__xnor2_2 _5739_ (.A(_1205_),
    .B(_1206_),
    .Y(_1207_));
 sky130_fd_sc_hd__and3_1 _5740_ (.A(_3423_),
    .B(_2248_),
    .C(_3573_),
    .X(_1208_));
 sky130_fd_sc_hd__a31o_1 _5741_ (.A1(_2160_),
    .A2(_3620_),
    .A3(_1080_),
    .B1(_1208_),
    .X(_1210_));
 sky130_fd_sc_hd__xor2_1 _5742_ (.A(_1207_),
    .B(_1210_),
    .X(_1211_));
 sky130_fd_sc_hd__xor2_1 _5743_ (.A(_1202_),
    .B(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__o21a_2 _5744_ (.A1(_1195_),
    .A2(_1196_),
    .B1(_1212_),
    .X(_1213_));
 sky130_fd_sc_hd__nor3_2 _5745_ (.A(_1195_),
    .B(_1196_),
    .C(_1212_),
    .Y(_1214_));
 sky130_fd_sc_hd__a211oi_4 _5746_ (.A1(_1193_),
    .A2(_1194_),
    .B1(_1213_),
    .C1(_1214_),
    .Y(_1215_));
 sky130_fd_sc_hd__o211a_1 _5747_ (.A1(_1213_),
    .A2(_1214_),
    .B1(_1193_),
    .C1(_1194_),
    .X(_1216_));
 sky130_fd_sc_hd__a41o_1 _5748_ (.A1(_3197_),
    .A2(_3272_),
    .A3(_2707_),
    .A4(_2751_),
    .B1(_1097_),
    .X(_1217_));
 sky130_fd_sc_hd__a32o_1 _5749_ (.A1(_0042_),
    .A2(_2773_),
    .A3(_1103_),
    .B1(_1102_),
    .B2(_2532_),
    .X(_1218_));
 sky130_fd_sc_hd__and4_1 _5750_ (.A(_3433_),
    .B(_3270_),
    .C(net6),
    .D(net7),
    .X(_1219_));
 sky130_fd_sc_hd__a22oi_1 _5751_ (.A1(_3633_),
    .A2(net6),
    .B1(_0380_),
    .B2(_3195_),
    .Y(_1221_));
 sky130_fd_sc_hd__and4bb_1 _5752_ (.A_N(_1219_),
    .B_N(_1221_),
    .C(_3343_),
    .D(_2686_),
    .X(_1222_));
 sky130_fd_sc_hd__o2bb2a_1 _5753_ (.A1_N(_3430_),
    .A2_N(_2696_),
    .B1(_1219_),
    .B2(_1221_),
    .X(_1223_));
 sky130_fd_sc_hd__or2_1 _5754_ (.A(_1222_),
    .B(_1223_),
    .X(_1224_));
 sky130_fd_sc_hd__xnor2_1 _5755_ (.A(_1218_),
    .B(_1224_),
    .Y(_1225_));
 sky130_fd_sc_hd__xnor2_1 _5756_ (.A(_1217_),
    .B(_1225_),
    .Y(_1226_));
 sky130_fd_sc_hd__and3_1 _5757_ (.A(_3352_),
    .B(_0373_),
    .C(net9),
    .X(_1227_));
 sky130_fd_sc_hd__a22o_1 _5758_ (.A1(_0373_),
    .A2(net9),
    .B1(net10),
    .B2(_3352_),
    .X(_1228_));
 sky130_fd_sc_hd__a21bo_1 _5759_ (.A1(_2565_),
    .A2(_1227_),
    .B1_N(_1228_),
    .X(_1229_));
 sky130_fd_sc_hd__nand2_1 _5760_ (.A(_0042_),
    .B(_2499_),
    .Y(_1230_));
 sky130_fd_sc_hd__xor2_1 _5761_ (.A(_1229_),
    .B(_1230_),
    .X(_1232_));
 sky130_fd_sc_hd__and2_1 _5762_ (.A(_0292_),
    .B(net11),
    .X(_1233_));
 sky130_fd_sc_hd__nand4_2 _5763_ (.A(_3451_),
    .B(_3452_),
    .C(_1854_),
    .D(_1887_),
    .Y(_1234_));
 sky130_fd_sc_hd__a22o_1 _5764_ (.A1(_0390_),
    .A2(net13),
    .B1(_1887_),
    .B2(_0488_),
    .X(_1235_));
 sky130_fd_sc_hd__nand3_1 _5765_ (.A(_1233_),
    .B(_1234_),
    .C(_1235_),
    .Y(_1236_));
 sky130_fd_sc_hd__a21o_1 _5766_ (.A1(_1234_),
    .A2(_1235_),
    .B1(_1233_),
    .X(_1237_));
 sky130_fd_sc_hd__a21bo_1 _5767_ (.A1(_1107_),
    .A2(_1109_),
    .B1_N(_1108_),
    .X(_1238_));
 sky130_fd_sc_hd__nand3_1 _5768_ (.A(_1236_),
    .B(_1237_),
    .C(_1238_),
    .Y(_1239_));
 sky130_fd_sc_hd__a21o_1 _5769_ (.A1(_1236_),
    .A2(_1237_),
    .B1(_1238_),
    .X(_1240_));
 sky130_fd_sc_hd__nand3_1 _5770_ (.A(_1232_),
    .B(_1239_),
    .C(_1240_),
    .Y(_1241_));
 sky130_fd_sc_hd__a21o_1 _5771_ (.A1(_1239_),
    .A2(_1240_),
    .B1(_1232_),
    .X(_1243_));
 sky130_fd_sc_hd__a21bo_1 _5772_ (.A1(_1106_),
    .A2(_1115_),
    .B1_N(_1114_),
    .X(_1244_));
 sky130_fd_sc_hd__and3_2 _5773_ (.A(_1241_),
    .B(_1243_),
    .C(_1244_),
    .X(_1245_));
 sky130_fd_sc_hd__a21oi_2 _5774_ (.A1(_1241_),
    .A2(_1243_),
    .B1(_1244_),
    .Y(_1246_));
 sky130_fd_sc_hd__or3_2 _5775_ (.A(_1226_),
    .B(_1245_),
    .C(_1246_),
    .X(_1247_));
 sky130_fd_sc_hd__o21ai_2 _5776_ (.A1(_1245_),
    .A2(_1246_),
    .B1(_1226_),
    .Y(_1248_));
 sky130_fd_sc_hd__o211ai_4 _5777_ (.A1(_1119_),
    .A2(net128),
    .B1(_1247_),
    .C1(_1248_),
    .Y(_1249_));
 sky130_fd_sc_hd__a211o_1 _5778_ (.A1(_1247_),
    .A2(_1248_),
    .B1(_1119_),
    .C1(_1121_),
    .X(_1250_));
 sky130_fd_sc_hd__and4bb_1 _5779_ (.A_N(_1215_),
    .B_N(_1216_),
    .C(_1249_),
    .D(_1250_),
    .X(_1251_));
 sky130_fd_sc_hd__a2bb2oi_2 _5780_ (.A1_N(_1215_),
    .A2_N(_1216_),
    .B1(_1249_),
    .B2(_1250_),
    .Y(_1252_));
 sky130_fd_sc_hd__a211oi_4 _5781_ (.A1(_1124_),
    .A2(net137),
    .B1(_1251_),
    .C1(_1252_),
    .Y(_1254_));
 sky130_fd_sc_hd__o211a_1 _5782_ (.A1(_1251_),
    .A2(_1252_),
    .B1(_1124_),
    .C1(net137),
    .X(_1255_));
 sky130_fd_sc_hd__or4_2 _5783_ (.A(net107),
    .B(_1192_),
    .C(_1254_),
    .D(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__o22ai_4 _5784_ (.A1(net107),
    .A2(_1192_),
    .B1(_1254_),
    .B2(_1255_),
    .Y(_1257_));
 sky130_fd_sc_hd__o211ai_2 _5785_ (.A1(_1128_),
    .A2(net199),
    .B1(_1256_),
    .C1(_1257_),
    .Y(_1258_));
 sky130_fd_sc_hd__a211o_1 _5786_ (.A1(_1256_),
    .A2(_1257_),
    .B1(_1128_),
    .C1(_1158_),
    .X(_1259_));
 sky130_fd_sc_hd__and3_1 _5787_ (.A(_1157_),
    .B(_1258_),
    .C(_1259_),
    .X(_1260_));
 sky130_fd_sc_hd__a21oi_1 _5788_ (.A1(_1258_),
    .A2(_1259_),
    .B1(_1157_),
    .Y(_1261_));
 sky130_fd_sc_hd__nor2_2 _5789_ (.A(_1260_),
    .B(_1261_),
    .Y(_1262_));
 sky130_fd_sc_hd__or2b_2 _5790_ (.A(_1132_),
    .B_N(_1135_),
    .X(_1263_));
 sky130_fd_sc_hd__xnor2_2 _5791_ (.A(_1262_),
    .B(_1263_),
    .Y(_1265_));
 sky130_fd_sc_hd__a21bo_1 _5792_ (.A1(net132),
    .A2(_1139_),
    .B1_N(_1138_),
    .X(_1266_));
 sky130_fd_sc_hd__xor2_2 _5793_ (.A(_1265_),
    .B(_1266_),
    .X(_1267_));
 sky130_fd_sc_hd__a21oi_1 _5794_ (.A1(_1151_),
    .A2(_1155_),
    .B1(_1267_),
    .Y(_1268_));
 sky130_fd_sc_hd__a31o_1 _5795_ (.A1(_1151_),
    .A2(_1267_),
    .A3(_1155_),
    .B1(_3192_),
    .X(_1269_));
 sky130_fd_sc_hd__or2_2 _5796_ (.A(_1909_),
    .B(_1170_),
    .X(_1270_));
 sky130_fd_sc_hd__nand2_2 _5797_ (.A(_1909_),
    .B(_1170_),
    .Y(_1271_));
 sky130_fd_sc_hd__nand2_4 _5798_ (.A(_1270_),
    .B(_1271_),
    .Y(_1272_));
 sky130_fd_sc_hd__and2b_1 _5799_ (.A_N(_1008_),
    .B(_1876_),
    .X(_1273_));
 sky130_fd_sc_hd__a21o_1 _5800_ (.A1(_1011_),
    .A2(_1014_),
    .B1(_1273_),
    .X(_1274_));
 sky130_fd_sc_hd__xor2_1 _5801_ (.A(_1272_),
    .B(_1274_),
    .X(_1276_));
 sky130_fd_sc_hd__clkbuf_4 _5802_ (.A(_0000_),
    .X(_1277_));
 sky130_fd_sc_hd__a21o_1 _5803_ (.A1(_0438_),
    .A2(_1271_),
    .B1(_1277_),
    .X(_1278_));
 sky130_fd_sc_hd__o22ai_1 _5804_ (.A1(_3712_),
    .A2(_1270_),
    .B1(_1271_),
    .B2(_0309_),
    .Y(_1279_));
 sky130_fd_sc_hd__o21a_1 _5805_ (.A1(_0848_),
    .A2(_3200_),
    .B1(_3161_),
    .X(_1280_));
 sky130_fd_sc_hd__and3_1 _5806_ (.A(_0848_),
    .B(_3097_),
    .C(_3126_),
    .X(_1281_));
 sky130_fd_sc_hd__a2111o_1 _5807_ (.A1(_1270_),
    .A2(_1278_),
    .B1(_1279_),
    .C1(_1280_),
    .D1(_1281_),
    .X(_1282_));
 sky130_fd_sc_hd__mux4_1 _5808_ (.A0(_1909_),
    .A1(_1876_),
    .A2(_0862_),
    .A3(_2587_),
    .S0(_0583_),
    .S1(_0584_),
    .X(_1283_));
 sky130_fd_sc_hd__mux2_1 _5809_ (.A0(_0710_),
    .A1(_1283_),
    .S(_0429_),
    .X(_1284_));
 sky130_fd_sc_hd__mux2_1 _5810_ (.A0(_0188_),
    .A1(_1284_),
    .S(_0189_),
    .X(_1285_));
 sky130_fd_sc_hd__nand2_1 _5811_ (.A(_0844_),
    .B(_1285_),
    .Y(_1287_));
 sky130_fd_sc_hd__a21oi_1 _5812_ (.A1(_3155_),
    .A2(_1287_),
    .B1(_0861_),
    .Y(_1288_));
 sky130_fd_sc_hd__a21oi_1 _5813_ (.A1(_1021_),
    .A2(_1029_),
    .B1(_1272_),
    .Y(_1289_));
 sky130_fd_sc_hd__a31o_1 _5814_ (.A1(_1021_),
    .A2(_1029_),
    .A3(_1272_),
    .B1(_3596_),
    .X(_1290_));
 sky130_fd_sc_hd__or2_1 _5815_ (.A(_1289_),
    .B(_1290_),
    .X(_1291_));
 sky130_fd_sc_hd__or3b_2 _5816_ (.A(_1282_),
    .B(_1288_),
    .C_N(_1291_),
    .X(_1292_));
 sky130_fd_sc_hd__a21oi_4 _5817_ (.A1(_3571_),
    .A2(_1276_),
    .B1(_1292_),
    .Y(_1293_));
 sky130_fd_sc_hd__o21ai_4 _5818_ (.A1(_1268_),
    .A2(_1269_),
    .B1(_1293_),
    .Y(net82));
 sky130_fd_sc_hd__clkbuf_4 _5819_ (.A(net47),
    .X(_1294_));
 sky130_fd_sc_hd__clkbuf_4 _5820_ (.A(_1294_),
    .X(_1295_));
 sky130_fd_sc_hd__and2_1 _5821_ (.A(_1942_),
    .B(_1295_),
    .X(_1297_));
 sky130_fd_sc_hd__nor2_1 _5822_ (.A(_1942_),
    .B(_1295_),
    .Y(_1298_));
 sky130_fd_sc_hd__or2_2 _5823_ (.A(_1297_),
    .B(_1298_),
    .X(_1299_));
 sky130_fd_sc_hd__and2b_1 _5824_ (.A_N(_1170_),
    .B(_1909_),
    .X(_1300_));
 sky130_fd_sc_hd__a21o_1 _5825_ (.A1(_1272_),
    .A2(_1274_),
    .B1(_1300_),
    .X(_1301_));
 sky130_fd_sc_hd__or2_1 _5826_ (.A(_1299_),
    .B(_1301_),
    .X(_1302_));
 sky130_fd_sc_hd__nand2_1 _5827_ (.A(_1299_),
    .B(_1301_),
    .Y(_1303_));
 sky130_fd_sc_hd__nand2_1 _5828_ (.A(_1010_),
    .B(_1270_),
    .Y(_1304_));
 sky130_fd_sc_hd__o311ai_4 _5829_ (.A1(_1011_),
    .A2(_1027_),
    .A3(_1272_),
    .B1(_1304_),
    .C1(_1271_),
    .Y(_1305_));
 sky130_fd_sc_hd__xnor2_1 _5830_ (.A(_1299_),
    .B(_1305_),
    .Y(_1306_));
 sky130_fd_sc_hd__mux4_1 _5831_ (.A0(_1942_),
    .A1(_1909_),
    .A2(_1876_),
    .A3(_0862_),
    .S0(_0583_),
    .S1(_0864_),
    .X(_1308_));
 sky130_fd_sc_hd__mux2_1 _5832_ (.A0(_0845_),
    .A1(_1308_),
    .S(_0866_),
    .X(_1309_));
 sky130_fd_sc_hd__mux2_1 _5833_ (.A0(_0305_),
    .A1(_1309_),
    .S(_0867_),
    .X(_1310_));
 sky130_fd_sc_hd__a21bo_1 _5834_ (.A1(_0844_),
    .A2(_1310_),
    .B1_N(_3228_),
    .X(_1311_));
 sky130_fd_sc_hd__o21ba_1 _5835_ (.A1(_3589_),
    .A2(_1297_),
    .B1_N(_1277_),
    .X(_1312_));
 sky130_fd_sc_hd__nor2_1 _5836_ (.A(_1298_),
    .B(_1312_),
    .Y(_1313_));
 sky130_fd_sc_hd__a221o_1 _5837_ (.A1(_0854_),
    .A2(_1297_),
    .B1(_1298_),
    .B2(_0855_),
    .C1(_1280_),
    .X(_1314_));
 sky130_fd_sc_hd__a311o_1 _5838_ (.A1(_0861_),
    .A2(_3126_),
    .A3(_3213_),
    .B1(_1313_),
    .C1(_1314_),
    .X(_1315_));
 sky130_fd_sc_hd__a221o_1 _5839_ (.A1(_0419_),
    .A2(_1306_),
    .B1(_1311_),
    .B2(_0573_),
    .C1(_1315_),
    .X(_1316_));
 sky130_fd_sc_hd__or3_1 _5840_ (.A(_0904_),
    .B(_1043_),
    .C(_1156_),
    .X(_1317_));
 sky130_fd_sc_hd__inv_2 _5841_ (.A(_1317_),
    .Y(_1319_));
 sky130_fd_sc_hd__nor2_1 _5842_ (.A(_1189_),
    .B(_1191_),
    .Y(_1320_));
 sky130_fd_sc_hd__and2b_1 _5843_ (.A_N(_1166_),
    .B(_1167_),
    .X(_1321_));
 sky130_fd_sc_hd__a31oi_4 _5844_ (.A1(_3209_),
    .A2(_1170_),
    .A3(_1168_),
    .B1(_1321_),
    .Y(_1322_));
 sky130_fd_sc_hd__xnor2_1 _5845_ (.A(_1320_),
    .B(_1322_),
    .Y(_1323_));
 sky130_fd_sc_hd__nor4_1 _5846_ (.A(_1191_),
    .B(_1192_),
    .C(_1254_),
    .D(_1255_),
    .Y(_1324_));
 sky130_fd_sc_hd__a22o_1 _5847_ (.A1(_0434_),
    .A2(net46),
    .B1(_1294_),
    .B2(_0466_),
    .X(_1325_));
 sky130_fd_sc_hd__inv_2 _5848_ (.A(_1325_),
    .Y(_1326_));
 sky130_fd_sc_hd__and4_1 _5849_ (.A(_0707_),
    .B(_0477_),
    .C(_1169_),
    .D(_1294_),
    .X(_1327_));
 sky130_fd_sc_hd__or2_1 _5850_ (.A(_1326_),
    .B(_1327_),
    .X(_1328_));
 sky130_fd_sc_hd__and4_1 _5851_ (.A(_0085_),
    .B(_1264_),
    .C(net42),
    .D(net43),
    .X(_1330_));
 sky130_fd_sc_hd__inv_2 _5852_ (.A(_1330_),
    .Y(_1331_));
 sky130_fd_sc_hd__a22o_1 _5853_ (.A1(_3440_),
    .A2(_0720_),
    .B1(_0873_),
    .B2(_1275_),
    .X(_1332_));
 sky130_fd_sc_hd__and4_1 _5854_ (.A(_0335_),
    .B(net45),
    .C(_1331_),
    .D(_1332_),
    .X(_1333_));
 sky130_fd_sc_hd__a22oi_1 _5855_ (.A1(_0346_),
    .A2(net45),
    .B1(_1331_),
    .B2(_1332_),
    .Y(_1334_));
 sky130_fd_sc_hd__or2_2 _5856_ (.A(_1333_),
    .B(_1334_),
    .X(_1335_));
 sky130_fd_sc_hd__or2_2 _5857_ (.A(_1160_),
    .B(_1163_),
    .X(_1336_));
 sky130_fd_sc_hd__xor2_4 _5858_ (.A(_1335_),
    .B(_1336_),
    .X(_1337_));
 sky130_fd_sc_hd__xnor2_2 _5859_ (.A(_1328_),
    .B(_1337_),
    .Y(_1338_));
 sky130_fd_sc_hd__nand2_1 _5860_ (.A(_1174_),
    .B(_1182_),
    .Y(_1339_));
 sky130_fd_sc_hd__or2_1 _5861_ (.A(_1175_),
    .B(_1178_),
    .X(_1341_));
 sky130_fd_sc_hd__and4_1 _5862_ (.A(_2368_),
    .B(_2423_),
    .C(_0325_),
    .D(_0452_),
    .X(_1342_));
 sky130_fd_sc_hd__a22oi_1 _5863_ (.A1(_2434_),
    .A2(_0325_),
    .B1(_0452_),
    .B2(_3442_),
    .Y(_1343_));
 sky130_fd_sc_hd__and4bb_1 _5864_ (.A_N(_1342_),
    .B_N(_1343_),
    .C(_2313_),
    .D(net41),
    .X(_1344_));
 sky130_fd_sc_hd__o2bb2a_1 _5865_ (.A1_N(_2313_),
    .A2_N(_0654_),
    .B1(_1342_),
    .B2(_1343_),
    .X(_1345_));
 sky130_fd_sc_hd__a211o_1 _5866_ (.A1(_1197_),
    .A2(_1200_),
    .B1(_1344_),
    .C1(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__o211ai_1 _5867_ (.A1(_1344_),
    .A2(_1345_),
    .B1(_1197_),
    .C1(_1200_),
    .Y(_1347_));
 sky130_fd_sc_hd__and2_1 _5868_ (.A(_1346_),
    .B(_1347_),
    .X(_1348_));
 sky130_fd_sc_hd__xnor2_2 _5869_ (.A(_1341_),
    .B(_1348_),
    .Y(_1349_));
 sky130_fd_sc_hd__a21oi_4 _5870_ (.A1(_1180_),
    .A2(_1339_),
    .B1(_1349_),
    .Y(_1350_));
 sky130_fd_sc_hd__and3_1 _5871_ (.A(_1180_),
    .B(_1339_),
    .C(_1349_),
    .X(_1352_));
 sky130_fd_sc_hd__or3_1 _5872_ (.A(_1338_),
    .B(_1350_),
    .C(_1352_),
    .X(_1353_));
 sky130_fd_sc_hd__o21ai_1 _5873_ (.A1(_1350_),
    .A2(_1352_),
    .B1(_1338_),
    .Y(_1354_));
 sky130_fd_sc_hd__o211a_1 _5874_ (.A1(_1213_),
    .A2(_1215_),
    .B1(_1353_),
    .C1(_1354_),
    .X(_1355_));
 sky130_fd_sc_hd__a211oi_2 _5875_ (.A1(_1353_),
    .A2(_1354_),
    .B1(_1213_),
    .C1(_1215_),
    .Y(_1356_));
 sky130_fd_sc_hd__a211oi_2 _5876_ (.A1(_1184_),
    .A2(_1186_),
    .B1(_1355_),
    .C1(_1356_),
    .Y(_1357_));
 sky130_fd_sc_hd__o211a_1 _5877_ (.A1(_1355_),
    .A2(_1356_),
    .B1(_1184_),
    .C1(_1186_),
    .X(_1358_));
 sky130_fd_sc_hd__or4bb_1 _5878_ (.A(_1215_),
    .B(_1216_),
    .C_N(_1249_),
    .D_N(_1250_),
    .X(_1359_));
 sky130_fd_sc_hd__or2b_1 _5879_ (.A(_1207_),
    .B_N(_1210_),
    .X(_1360_));
 sky130_fd_sc_hd__or2_1 _5880_ (.A(_1202_),
    .B(_1211_),
    .X(_1361_));
 sky130_fd_sc_hd__and2b_1 _5881_ (.A_N(_1224_),
    .B(_1218_),
    .X(_1363_));
 sky130_fd_sc_hd__and2_1 _5882_ (.A(_1217_),
    .B(_1225_),
    .X(_1364_));
 sky130_fd_sc_hd__and4_1 _5883_ (.A(_0247_),
    .B(_2204_),
    .C(_3718_),
    .D(_0099_),
    .X(_1365_));
 sky130_fd_sc_hd__a22o_1 _5884_ (.A1(_2204_),
    .A2(_3718_),
    .B1(_0099_),
    .B2(_0247_),
    .X(_1366_));
 sky130_fd_sc_hd__or2b_1 _5885_ (.A(_1365_),
    .B_N(_1366_),
    .X(_1367_));
 sky130_fd_sc_hd__nand2_1 _5886_ (.A(_2117_),
    .B(_0220_),
    .Y(_1368_));
 sky130_fd_sc_hd__xnor2_2 _5887_ (.A(_1367_),
    .B(_1368_),
    .Y(_1369_));
 sky130_fd_sc_hd__nand4_1 _5888_ (.A(_3423_),
    .B(_0105_),
    .C(_0491_),
    .D(_2696_),
    .Y(_1370_));
 sky130_fd_sc_hd__a22o_1 _5889_ (.A1(_3511_),
    .A2(_0491_),
    .B1(_2686_),
    .B2(_0104_),
    .X(_1371_));
 sky130_fd_sc_hd__and3_1 _5890_ (.A(_3709_),
    .B(_1370_),
    .C(_1371_),
    .X(_1372_));
 sky130_fd_sc_hd__a21oi_1 _5891_ (.A1(_1370_),
    .A2(_1371_),
    .B1(_3709_),
    .Y(_1374_));
 sky130_fd_sc_hd__nor2_1 _5892_ (.A(_1372_),
    .B(_1374_),
    .Y(_1375_));
 sky130_fd_sc_hd__a31o_1 _5893_ (.A1(_2215_),
    .A2(_3620_),
    .A3(_1204_),
    .B1(_1203_),
    .X(_1376_));
 sky130_fd_sc_hd__xor2_2 _5894_ (.A(_1375_),
    .B(_1376_),
    .X(_1377_));
 sky130_fd_sc_hd__xnor2_2 _5895_ (.A(_1369_),
    .B(_1377_),
    .Y(_1378_));
 sky130_fd_sc_hd__o21a_2 _5896_ (.A1(_1363_),
    .A2(_1364_),
    .B1(_1378_),
    .X(_1379_));
 sky130_fd_sc_hd__nor3_2 _5897_ (.A(_1363_),
    .B(_1364_),
    .C(_1378_),
    .Y(_1380_));
 sky130_fd_sc_hd__a211oi_4 _5898_ (.A1(_1360_),
    .A2(_1361_),
    .B1(_1379_),
    .C1(_1380_),
    .Y(_1381_));
 sky130_fd_sc_hd__o211a_1 _5899_ (.A1(_1379_),
    .A2(_1380_),
    .B1(_1360_),
    .C1(_1361_),
    .X(_1382_));
 sky130_fd_sc_hd__nor3_1 _5900_ (.A(_1226_),
    .B(_1245_),
    .C(_1246_),
    .Y(_1383_));
 sky130_fd_sc_hd__or2_1 _5901_ (.A(_1219_),
    .B(_1222_),
    .X(_1385_));
 sky130_fd_sc_hd__a32o_1 _5902_ (.A1(_2881_),
    .A2(_2489_),
    .A3(_1228_),
    .B1(_1227_),
    .B2(_2565_),
    .X(_1386_));
 sky130_fd_sc_hd__nand4_2 _5903_ (.A(_3632_),
    .B(_3633_),
    .C(_0380_),
    .D(_2489_),
    .Y(_1387_));
 sky130_fd_sc_hd__a22o_1 _5904_ (.A1(_3633_),
    .A2(net7),
    .B1(net8),
    .B2(_3195_),
    .X(_1388_));
 sky130_fd_sc_hd__nand4_1 _5905_ (.A(_3631_),
    .B(_2751_),
    .C(_1387_),
    .D(_1388_),
    .Y(_1389_));
 sky130_fd_sc_hd__a22o_1 _5906_ (.A1(_3430_),
    .A2(_2740_),
    .B1(_1387_),
    .B2(_1388_),
    .X(_1390_));
 sky130_fd_sc_hd__and3_1 _5907_ (.A(_1386_),
    .B(_1389_),
    .C(_1390_),
    .X(_1391_));
 sky130_fd_sc_hd__a21o_1 _5908_ (.A1(_1389_),
    .A2(_1390_),
    .B1(_1386_),
    .X(_1392_));
 sky130_fd_sc_hd__and2b_1 _5909_ (.A_N(_1391_),
    .B(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__xnor2_1 _5910_ (.A(_1385_),
    .B(_1393_),
    .Y(_1394_));
 sky130_fd_sc_hd__and3_1 _5911_ (.A(_0161_),
    .B(_0373_),
    .C(_2565_),
    .X(_1396_));
 sky130_fd_sc_hd__a22o_1 _5912_ (.A1(_3531_),
    .A2(net10),
    .B1(net11),
    .B2(_0161_),
    .X(_1397_));
 sky130_fd_sc_hd__a21bo_1 _5913_ (.A1(_2598_),
    .A2(_1396_),
    .B1_N(_1397_),
    .X(_1398_));
 sky130_fd_sc_hd__nand2_1 _5914_ (.A(_0042_),
    .B(_2532_),
    .Y(_1399_));
 sky130_fd_sc_hd__xor2_1 _5915_ (.A(_1398_),
    .B(_1399_),
    .X(_1400_));
 sky130_fd_sc_hd__nand4_1 _5916_ (.A(_0488_),
    .B(_0390_),
    .C(_1887_),
    .D(net15),
    .Y(_1401_));
 sky130_fd_sc_hd__a22o_1 _5917_ (.A1(net178),
    .A2(_1887_),
    .B1(net15),
    .B2(_3242_),
    .X(_1402_));
 sky130_fd_sc_hd__and2_1 _5918_ (.A(_0281_),
    .B(net13),
    .X(_1403_));
 sky130_fd_sc_hd__nand3_1 _5919_ (.A(_1401_),
    .B(_1402_),
    .C(_1403_),
    .Y(_1404_));
 sky130_fd_sc_hd__a21o_1 _5920_ (.A1(_1401_),
    .A2(_1402_),
    .B1(_1403_),
    .X(_1405_));
 sky130_fd_sc_hd__a21bo_1 _5921_ (.A1(_1233_),
    .A2(_1235_),
    .B1_N(_1234_),
    .X(_1407_));
 sky130_fd_sc_hd__nand3_1 _5922_ (.A(_1404_),
    .B(_1405_),
    .C(_1407_),
    .Y(_1408_));
 sky130_fd_sc_hd__a21o_1 _5923_ (.A1(_1404_),
    .A2(_1405_),
    .B1(_1407_),
    .X(_1409_));
 sky130_fd_sc_hd__nand3_1 _5924_ (.A(_1400_),
    .B(_1408_),
    .C(_1409_),
    .Y(_1410_));
 sky130_fd_sc_hd__a21o_1 _5925_ (.A1(_1408_),
    .A2(_1409_),
    .B1(_1400_),
    .X(_1411_));
 sky130_fd_sc_hd__a21bo_1 _5926_ (.A1(_1232_),
    .A2(_1240_),
    .B1_N(_1239_),
    .X(_1412_));
 sky130_fd_sc_hd__and3_2 _5927_ (.A(_1410_),
    .B(_1411_),
    .C(_1412_),
    .X(_1413_));
 sky130_fd_sc_hd__a21oi_2 _5928_ (.A1(_1410_),
    .A2(_1411_),
    .B1(_1412_),
    .Y(_1414_));
 sky130_fd_sc_hd__or3_1 _5929_ (.A(_1394_),
    .B(_1413_),
    .C(_1414_),
    .X(_1415_));
 sky130_fd_sc_hd__o21ai_1 _5930_ (.A1(_1413_),
    .A2(_1414_),
    .B1(_1394_),
    .Y(_1416_));
 sky130_fd_sc_hd__o211a_2 _5931_ (.A1(_1245_),
    .A2(_1383_),
    .B1(_1415_),
    .C1(_1416_),
    .X(_1418_));
 sky130_fd_sc_hd__a211oi_2 _5932_ (.A1(_1415_),
    .A2(_1416_),
    .B1(_1245_),
    .C1(_1383_),
    .Y(_1419_));
 sky130_fd_sc_hd__nor4_1 _5933_ (.A(_1381_),
    .B(_1382_),
    .C(_1418_),
    .D(_1419_),
    .Y(_1420_));
 sky130_fd_sc_hd__o22a_1 _5934_ (.A1(_1381_),
    .A2(_1382_),
    .B1(_1418_),
    .B2(_1419_),
    .X(_1421_));
 sky130_fd_sc_hd__a211o_1 _5935_ (.A1(_1249_),
    .A2(_1359_),
    .B1(net203),
    .C1(_1421_),
    .X(_1422_));
 sky130_fd_sc_hd__o211ai_1 _5936_ (.A1(net203),
    .A2(_1421_),
    .B1(_1249_),
    .C1(_1359_),
    .Y(_1423_));
 sky130_fd_sc_hd__or4bb_2 _5937_ (.A(_1357_),
    .B(_1358_),
    .C_N(_1422_),
    .D_N(_1423_),
    .X(_1424_));
 sky130_fd_sc_hd__a2bb2o_1 _5938_ (.A1_N(_1357_),
    .A2_N(_1358_),
    .B1(_1422_),
    .B2(_1423_),
    .X(_1425_));
 sky130_fd_sc_hd__o211a_1 _5939_ (.A1(_1254_),
    .A2(_1324_),
    .B1(_1424_),
    .C1(_1425_),
    .X(_1426_));
 sky130_fd_sc_hd__a211oi_2 _5940_ (.A1(_1424_),
    .A2(_1425_),
    .B1(_1254_),
    .C1(net198),
    .Y(_1427_));
 sky130_fd_sc_hd__or3_1 _5941_ (.A(_1323_),
    .B(_1426_),
    .C(_1427_),
    .X(_1429_));
 sky130_fd_sc_hd__o21ai_1 _5942_ (.A1(_1426_),
    .A2(_1427_),
    .B1(_1323_),
    .Y(_1430_));
 sky130_fd_sc_hd__nand2_2 _5943_ (.A(_1429_),
    .B(_1430_),
    .Y(_1431_));
 sky130_fd_sc_hd__a21bo_2 _5944_ (.A1(_1157_),
    .A2(_1259_),
    .B1_N(_1258_),
    .X(_1432_));
 sky130_fd_sc_hd__xnor2_4 _5945_ (.A(_1431_),
    .B(_1432_),
    .Y(_1433_));
 sky130_fd_sc_hd__xnor2_4 _5946_ (.A(_1319_),
    .B(_1433_),
    .Y(_1434_));
 sky130_fd_sc_hd__nand2_1 _5947_ (.A(_1262_),
    .B(_1263_),
    .Y(_1435_));
 sky130_fd_sc_hd__o21a_1 _5948_ (.A1(_1138_),
    .A2(_1265_),
    .B1(_1435_),
    .X(_1436_));
 sky130_fd_sc_hd__xnor2_2 _5949_ (.A(_1434_),
    .B(_1436_),
    .Y(_1437_));
 sky130_fd_sc_hd__nand3_1 _5950_ (.A(net133),
    .B(_1138_),
    .C(_1139_),
    .Y(_1438_));
 sky130_fd_sc_hd__o22a_1 _5951_ (.A1(_1265_),
    .A2(_1438_),
    .B1(_1267_),
    .B2(_1155_),
    .X(_1440_));
 sky130_fd_sc_hd__or2_1 _5952_ (.A(_1142_),
    .B(_1267_),
    .X(_1441_));
 sky130_fd_sc_hd__a21o_1 _5953_ (.A1(_1146_),
    .A2(_1149_),
    .B1(_1441_),
    .X(_1442_));
 sky130_fd_sc_hd__nand3_1 _5954_ (.A(_1437_),
    .B(_1440_),
    .C(_1442_),
    .Y(_1443_));
 sky130_fd_sc_hd__a21o_1 _5955_ (.A1(_1440_),
    .A2(_1442_),
    .B1(_1437_),
    .X(_1444_));
 sky130_fd_sc_hd__and3_1 _5956_ (.A(_0320_),
    .B(_1443_),
    .C(_1444_),
    .X(_1445_));
 sky130_fd_sc_hd__a311o_4 _5957_ (.A1(_3571_),
    .A2(_1302_),
    .A3(_1303_),
    .B1(_1316_),
    .C1(_1445_),
    .X(net83));
 sky130_fd_sc_hd__and2b_1 _5958_ (.A_N(_1295_),
    .B(_1942_),
    .X(_1446_));
 sky130_fd_sc_hd__inv_2 _5959_ (.A(_1446_),
    .Y(_1447_));
 sky130_fd_sc_hd__clkbuf_4 _5960_ (.A(net48),
    .X(_1448_));
 sky130_fd_sc_hd__or2_2 _5961_ (.A(_1963_),
    .B(_1448_),
    .X(_1450_));
 sky130_fd_sc_hd__nand2_2 _5962_ (.A(_1963_),
    .B(_1448_),
    .Y(_1451_));
 sky130_fd_sc_hd__and2_1 _5963_ (.A(_1450_),
    .B(_1451_),
    .X(_1452_));
 sky130_fd_sc_hd__a21o_1 _5964_ (.A1(_1303_),
    .A2(_1447_),
    .B1(_1452_),
    .X(_1453_));
 sky130_fd_sc_hd__nand2_1 _5965_ (.A(_1450_),
    .B(_1451_),
    .Y(_1454_));
 sky130_fd_sc_hd__or3b_1 _5966_ (.A(_1454_),
    .B(_1446_),
    .C_N(_1303_),
    .X(_1455_));
 sky130_fd_sc_hd__nor2_1 _5967_ (.A(_1297_),
    .B(_1298_),
    .Y(_1456_));
 sky130_fd_sc_hd__a21o_1 _5968_ (.A1(_1456_),
    .A2(_1305_),
    .B1(_1297_),
    .X(_1457_));
 sky130_fd_sc_hd__nand2_1 _5969_ (.A(_1452_),
    .B(_1457_),
    .Y(_1458_));
 sky130_fd_sc_hd__o21a_1 _5970_ (.A1(_1452_),
    .A2(_1457_),
    .B1(_0419_),
    .X(_1459_));
 sky130_fd_sc_hd__a21o_1 _5971_ (.A1(_3126_),
    .A2(_3285_),
    .B1(_3161_),
    .X(_1461_));
 sky130_fd_sc_hd__a21o_1 _5972_ (.A1(_0438_),
    .A2(_1451_),
    .B1(_1277_),
    .X(_1462_));
 sky130_fd_sc_hd__o31a_1 _5973_ (.A1(_3490_),
    .A2(_0863_),
    .A3(_0864_),
    .B1(_0199_),
    .X(_1463_));
 sky130_fd_sc_hd__o22ai_1 _5974_ (.A1(_3712_),
    .A2(_1450_),
    .B1(_1451_),
    .B2(_0309_),
    .Y(_1464_));
 sky130_fd_sc_hd__a221o_1 _5975_ (.A1(_1450_),
    .A2(_1462_),
    .B1(_1463_),
    .B2(_3161_),
    .C1(_1464_),
    .X(_1465_));
 sky130_fd_sc_hd__mux4_1 _5976_ (.A0(_1963_),
    .A1(_1942_),
    .A2(_1909_),
    .A3(_1876_),
    .S0(_0863_),
    .S1(_0864_),
    .X(_1466_));
 sky130_fd_sc_hd__mux2_1 _5977_ (.A0(_0865_),
    .A1(_1466_),
    .S(_0866_),
    .X(_1467_));
 sky130_fd_sc_hd__mux2_1 _5978_ (.A0(_0435_),
    .A1(_1467_),
    .S(_0867_),
    .X(_1468_));
 sky130_fd_sc_hd__nand2_1 _5979_ (.A(_0844_),
    .B(_1468_),
    .Y(_1469_));
 sky130_fd_sc_hd__a21oi_1 _5980_ (.A1(_3295_),
    .A2(_1469_),
    .B1(_0861_),
    .Y(_1470_));
 sky130_fd_sc_hd__a211o_1 _5981_ (.A1(_0861_),
    .A2(_1461_),
    .B1(_1465_),
    .C1(_1470_),
    .X(_1472_));
 sky130_fd_sc_hd__nor2_2 _5982_ (.A(_1320_),
    .B(_1322_),
    .Y(_1473_));
 sky130_fd_sc_hd__and2b_1 _5983_ (.A_N(_1335_),
    .B(_1336_),
    .X(_1474_));
 sky130_fd_sc_hd__and2_2 _5984_ (.A(_1327_),
    .B(_1474_),
    .X(_1475_));
 sky130_fd_sc_hd__nor2_1 _5985_ (.A(_1327_),
    .B(_1474_),
    .Y(_1476_));
 sky130_fd_sc_hd__o32ai_4 _5986_ (.A1(_1326_),
    .A2(_1327_),
    .A3(_1337_),
    .B1(_1475_),
    .B2(_1476_),
    .Y(_1477_));
 sky130_fd_sc_hd__o21ai_1 _5987_ (.A1(_1355_),
    .A2(_1357_),
    .B1(_1477_),
    .Y(_1478_));
 sky130_fd_sc_hd__or3_1 _5988_ (.A(_1355_),
    .B(_1357_),
    .C(_1477_),
    .X(_1479_));
 sky130_fd_sc_hd__and2_1 _5989_ (.A(_1478_),
    .B(_1479_),
    .X(_1480_));
 sky130_fd_sc_hd__nor3_2 _5990_ (.A(_1338_),
    .B(_1350_),
    .C(_1352_),
    .Y(_1481_));
 sky130_fd_sc_hd__and4_1 _5991_ (.A(_0346_),
    .B(_0707_),
    .C(net46),
    .D(_1294_),
    .X(_1483_));
 sky130_fd_sc_hd__a22o_1 _5992_ (.A1(_0335_),
    .A2(net46),
    .B1(net47),
    .B2(_0434_),
    .X(_1484_));
 sky130_fd_sc_hd__and4b_1 _5993_ (.A_N(_1483_),
    .B(_1484_),
    .C(_0991_),
    .D(net48),
    .X(_1485_));
 sky130_fd_sc_hd__inv_2 _5994_ (.A(_1484_),
    .Y(_1486_));
 sky130_fd_sc_hd__o2bb2a_1 _5995_ (.A1_N(_0991_),
    .A2_N(net48),
    .B1(_1483_),
    .B2(_1486_),
    .X(_1487_));
 sky130_fd_sc_hd__or2_1 _5996_ (.A(_1485_),
    .B(_1487_),
    .X(_1488_));
 sky130_fd_sc_hd__and4_1 _5997_ (.A(_0095_),
    .B(_2313_),
    .C(_0720_),
    .D(_0873_),
    .X(_1489_));
 sky130_fd_sc_hd__a22o_1 _5998_ (.A1(_2313_),
    .A2(_0720_),
    .B1(_0873_),
    .B2(_0095_),
    .X(_1490_));
 sky130_fd_sc_hd__and4b_1 _5999_ (.A_N(_1489_),
    .B(_1490_),
    .C(_0215_),
    .D(net45),
    .X(_1491_));
 sky130_fd_sc_hd__inv_2 _6000_ (.A(_1489_),
    .Y(_1492_));
 sky130_fd_sc_hd__a22oi_1 _6001_ (.A1(_0215_),
    .A2(_1007_),
    .B1(_1492_),
    .B2(_1490_),
    .Y(_1494_));
 sky130_fd_sc_hd__or2_1 _6002_ (.A(_1491_),
    .B(_1494_),
    .X(_1495_));
 sky130_fd_sc_hd__or2_2 _6003_ (.A(_1330_),
    .B(_1333_),
    .X(_1496_));
 sky130_fd_sc_hd__xor2_2 _6004_ (.A(_1495_),
    .B(_1496_),
    .X(_1497_));
 sky130_fd_sc_hd__xor2_2 _6005_ (.A(_1488_),
    .B(_1497_),
    .X(_1498_));
 sky130_fd_sc_hd__nand2_1 _6006_ (.A(_1341_),
    .B(_1348_),
    .Y(_1499_));
 sky130_fd_sc_hd__or2_1 _6007_ (.A(_1342_),
    .B(_1344_),
    .X(_1500_));
 sky130_fd_sc_hd__a31o_1 _6008_ (.A1(_2117_),
    .A2(_0219_),
    .A3(_1366_),
    .B1(_1365_),
    .X(_1501_));
 sky130_fd_sc_hd__nand4_2 _6009_ (.A(_3530_),
    .B(_2117_),
    .C(_0326_),
    .D(_0453_),
    .Y(_1502_));
 sky130_fd_sc_hd__a22o_1 _6010_ (.A1(_3644_),
    .A2(_0326_),
    .B1(_0453_),
    .B2(_3530_),
    .X(_1503_));
 sky130_fd_sc_hd__nand4_1 _6011_ (.A(_2390_),
    .B(_0688_),
    .C(_1502_),
    .D(_1503_),
    .Y(_1505_));
 sky130_fd_sc_hd__a22o_1 _6012_ (.A1(_2390_),
    .A2(_0654_),
    .B1(_1502_),
    .B2(_1503_),
    .X(_1506_));
 sky130_fd_sc_hd__and3_1 _6013_ (.A(_1501_),
    .B(_1505_),
    .C(_1506_),
    .X(_1507_));
 sky130_fd_sc_hd__a21o_1 _6014_ (.A1(_1505_),
    .A2(_1506_),
    .B1(_1501_),
    .X(_1508_));
 sky130_fd_sc_hd__and2b_1 _6015_ (.A_N(_1507_),
    .B(_1508_),
    .X(_1509_));
 sky130_fd_sc_hd__xnor2_1 _6016_ (.A(_1500_),
    .B(_1509_),
    .Y(_1510_));
 sky130_fd_sc_hd__a21o_1 _6017_ (.A1(_1346_),
    .A2(_1499_),
    .B1(_1510_),
    .X(_1511_));
 sky130_fd_sc_hd__nand3_1 _6018_ (.A(_1346_),
    .B(_1499_),
    .C(_1510_),
    .Y(_1512_));
 sky130_fd_sc_hd__nand3_2 _6019_ (.A(_1498_),
    .B(_1511_),
    .C(_1512_),
    .Y(_1513_));
 sky130_fd_sc_hd__a21o_1 _6020_ (.A1(_1511_),
    .A2(_1512_),
    .B1(_1498_),
    .X(_1514_));
 sky130_fd_sc_hd__o211ai_4 _6021_ (.A1(_1379_),
    .A2(_1381_),
    .B1(_1513_),
    .C1(_1514_),
    .Y(_1516_));
 sky130_fd_sc_hd__a211o_1 _6022_ (.A1(_1513_),
    .A2(_1514_),
    .B1(_1379_),
    .C1(_1381_),
    .X(_1517_));
 sky130_fd_sc_hd__o211ai_4 _6023_ (.A1(_1350_),
    .A2(_1481_),
    .B1(_1516_),
    .C1(_1517_),
    .Y(_1518_));
 sky130_fd_sc_hd__a211o_1 _6024_ (.A1(_1516_),
    .A2(_1517_),
    .B1(_1350_),
    .C1(_1481_),
    .X(_1519_));
 sky130_fd_sc_hd__nand2_1 _6025_ (.A(_1375_),
    .B(_1376_),
    .Y(_1520_));
 sky130_fd_sc_hd__or2b_1 _6026_ (.A(_1369_),
    .B_N(_1377_),
    .X(_1521_));
 sky130_fd_sc_hd__a21o_1 _6027_ (.A1(_1385_),
    .A2(_1392_),
    .B1(_1391_),
    .X(_1522_));
 sky130_fd_sc_hd__and3_1 _6028_ (.A(_2215_),
    .B(_2259_),
    .C(_0099_),
    .X(_1523_));
 sky130_fd_sc_hd__a22o_1 _6029_ (.A1(_2259_),
    .A2(_3718_),
    .B1(_0099_),
    .B2(_2204_),
    .X(_1524_));
 sky130_fd_sc_hd__a21bo_1 _6030_ (.A1(_3719_),
    .A2(_1523_),
    .B1_N(_1524_),
    .X(_1525_));
 sky130_fd_sc_hd__nand2_1 _6031_ (.A(_2160_),
    .B(_0220_),
    .Y(_1527_));
 sky130_fd_sc_hd__xor2_1 _6032_ (.A(_1525_),
    .B(_1527_),
    .X(_1528_));
 sky130_fd_sc_hd__and4_1 _6033_ (.A(_3424_),
    .B(_3512_),
    .C(_2653_),
    .D(_2707_),
    .X(_1529_));
 sky130_fd_sc_hd__nand4_4 _6034_ (.A(_3423_),
    .B(_0105_),
    .C(_2696_),
    .D(_2751_),
    .Y(_1530_));
 sky130_fd_sc_hd__a22o_1 _6035_ (.A1(_0105_),
    .A2(_2696_),
    .B1(_2740_),
    .B2(_0104_),
    .X(_1531_));
 sky130_fd_sc_hd__nand4_4 _6036_ (.A(_0110_),
    .B(_2653_),
    .C(_1530_),
    .D(_1531_),
    .Y(_1532_));
 sky130_fd_sc_hd__a22o_1 _6037_ (.A1(_3620_),
    .A2(_2653_),
    .B1(_1530_),
    .B2(_1531_),
    .X(_1533_));
 sky130_fd_sc_hd__o211ai_4 _6038_ (.A1(_1529_),
    .A2(_1372_),
    .B1(_1532_),
    .C1(_1533_),
    .Y(_1534_));
 sky130_fd_sc_hd__a211o_1 _6039_ (.A1(_1532_),
    .A2(_1533_),
    .B1(_1529_),
    .C1(_1372_),
    .X(_1535_));
 sky130_fd_sc_hd__nand3_2 _6040_ (.A(_1528_),
    .B(_1534_),
    .C(_1535_),
    .Y(_1536_));
 sky130_fd_sc_hd__a21o_1 _6041_ (.A1(_1534_),
    .A2(_1535_),
    .B1(_1528_),
    .X(_1538_));
 sky130_fd_sc_hd__and3_2 _6042_ (.A(_1522_),
    .B(_1536_),
    .C(_1538_),
    .X(_1539_));
 sky130_fd_sc_hd__a21oi_2 _6043_ (.A1(_1536_),
    .A2(_1538_),
    .B1(_1522_),
    .Y(_1540_));
 sky130_fd_sc_hd__a211oi_4 _6044_ (.A1(_1520_),
    .A2(_1521_),
    .B1(_1539_),
    .C1(_1540_),
    .Y(_1541_));
 sky130_fd_sc_hd__o211a_1 _6045_ (.A1(_1539_),
    .A2(_1540_),
    .B1(_1520_),
    .C1(_1521_),
    .X(_1542_));
 sky130_fd_sc_hd__nor3_1 _6046_ (.A(_1394_),
    .B(_1413_),
    .C(_1414_),
    .Y(_1543_));
 sky130_fd_sc_hd__nand2_1 _6047_ (.A(_1387_),
    .B(_1389_),
    .Y(_1544_));
 sky130_fd_sc_hd__a32o_1 _6048_ (.A1(_2881_),
    .A2(_2532_),
    .A3(_1397_),
    .B1(_1396_),
    .B2(_2598_),
    .X(_1545_));
 sky130_fd_sc_hd__nand4_2 _6049_ (.A(_3632_),
    .B(_3633_),
    .C(_2489_),
    .D(_2521_),
    .Y(_1546_));
 sky130_fd_sc_hd__a22o_1 _6050_ (.A1(_3633_),
    .A2(net8),
    .B1(_2521_),
    .B2(_3195_),
    .X(_1547_));
 sky130_fd_sc_hd__nand4_1 _6051_ (.A(_3631_),
    .B(_2773_),
    .C(_1546_),
    .D(_1547_),
    .Y(_1549_));
 sky130_fd_sc_hd__a22o_1 _6052_ (.A1(_3430_),
    .A2(_2773_),
    .B1(_1546_),
    .B2(_1547_),
    .X(_1550_));
 sky130_fd_sc_hd__and3_1 _6053_ (.A(_1545_),
    .B(_1549_),
    .C(_1550_),
    .X(_1551_));
 sky130_fd_sc_hd__a21o_1 _6054_ (.A1(_1549_),
    .A2(_1550_),
    .B1(_1545_),
    .X(_1552_));
 sky130_fd_sc_hd__and2b_1 _6055_ (.A_N(_1551_),
    .B(_1552_),
    .X(_1553_));
 sky130_fd_sc_hd__xnor2_2 _6056_ (.A(_1544_),
    .B(_1553_),
    .Y(_1554_));
 sky130_fd_sc_hd__nand4_1 _6057_ (.A(_0488_),
    .B(_0390_),
    .C(net15),
    .D(net16),
    .Y(_1555_));
 sky130_fd_sc_hd__a22o_1 _6058_ (.A1(net178),
    .A2(net15),
    .B1(net16),
    .B2(_3242_),
    .X(_1556_));
 sky130_fd_sc_hd__and2_1 _6059_ (.A(_0281_),
    .B(_1887_),
    .X(_1557_));
 sky130_fd_sc_hd__nand3_1 _6060_ (.A(_1555_),
    .B(_1556_),
    .C(_1557_),
    .Y(_1558_));
 sky130_fd_sc_hd__a21o_1 _6061_ (.A1(_1555_),
    .A2(_1556_),
    .B1(_1557_),
    .X(_1560_));
 sky130_fd_sc_hd__a21bo_1 _6062_ (.A1(_1402_),
    .A2(_1403_),
    .B1_N(_1401_),
    .X(_1561_));
 sky130_fd_sc_hd__nand3_1 _6063_ (.A(_1558_),
    .B(_1560_),
    .C(_1561_),
    .Y(_1562_));
 sky130_fd_sc_hd__a21o_1 _6064_ (.A1(_1558_),
    .A2(_1560_),
    .B1(_1561_),
    .X(_1563_));
 sky130_fd_sc_hd__and3_1 _6065_ (.A(_3169_),
    .B(net191),
    .C(net11),
    .X(_1564_));
 sky130_fd_sc_hd__a22o_1 _6066_ (.A1(_0030_),
    .A2(net11),
    .B1(net13),
    .B2(_3169_),
    .X(_1565_));
 sky130_fd_sc_hd__a21bo_1 _6067_ (.A1(_1854_),
    .A2(_1564_),
    .B1_N(_1565_),
    .X(_1566_));
 sky130_fd_sc_hd__nand2_1 _6068_ (.A(_2881_),
    .B(_2565_),
    .Y(_1567_));
 sky130_fd_sc_hd__xor2_1 _6069_ (.A(_1566_),
    .B(_1567_),
    .X(_1568_));
 sky130_fd_sc_hd__nand3_1 _6070_ (.A(_1562_),
    .B(_1563_),
    .C(_1568_),
    .Y(_1569_));
 sky130_fd_sc_hd__a21o_1 _6071_ (.A1(_1562_),
    .A2(_1563_),
    .B1(_1568_),
    .X(_1571_));
 sky130_fd_sc_hd__a21bo_1 _6072_ (.A1(_1400_),
    .A2(_1409_),
    .B1_N(_1408_),
    .X(_1572_));
 sky130_fd_sc_hd__and3_2 _6073_ (.A(_1569_),
    .B(_1571_),
    .C(_1572_),
    .X(_1573_));
 sky130_fd_sc_hd__a21oi_2 _6074_ (.A1(_1569_),
    .A2(_1571_),
    .B1(_1572_),
    .Y(_1574_));
 sky130_fd_sc_hd__or3_2 _6075_ (.A(_1554_),
    .B(_1573_),
    .C(_1574_),
    .X(_1575_));
 sky130_fd_sc_hd__o21ai_2 _6076_ (.A1(_1573_),
    .A2(_1574_),
    .B1(_1554_),
    .Y(_1576_));
 sky130_fd_sc_hd__o211ai_4 _6077_ (.A1(_1413_),
    .A2(net121),
    .B1(_1575_),
    .C1(_1576_),
    .Y(_1577_));
 sky130_fd_sc_hd__a211o_1 _6078_ (.A1(_1575_),
    .A2(_1576_),
    .B1(_1413_),
    .C1(_1543_),
    .X(_1578_));
 sky130_fd_sc_hd__or4bb_4 _6079_ (.A(_1541_),
    .B(_1542_),
    .C_N(_1577_),
    .D_N(_1578_),
    .X(_1579_));
 sky130_fd_sc_hd__a2bb2o_1 _6080_ (.A1_N(_1541_),
    .A2_N(_1542_),
    .B1(_1577_),
    .B2(_1578_),
    .X(_1580_));
 sky130_fd_sc_hd__o211ai_2 _6081_ (.A1(_1418_),
    .A2(net109),
    .B1(_1579_),
    .C1(_1580_),
    .Y(_1582_));
 sky130_fd_sc_hd__a211o_1 _6082_ (.A1(_1579_),
    .A2(_1580_),
    .B1(_1418_),
    .C1(net109),
    .X(_1583_));
 sky130_fd_sc_hd__and4_2 _6083_ (.A(_1518_),
    .B(_1519_),
    .C(_1582_),
    .D(_1583_),
    .X(_1584_));
 sky130_fd_sc_hd__a22oi_2 _6084_ (.A1(_1518_),
    .A2(_1519_),
    .B1(_1582_),
    .B2(_1583_),
    .Y(_1585_));
 sky130_fd_sc_hd__a211o_1 _6085_ (.A1(net154),
    .A2(_1424_),
    .B1(_1584_),
    .C1(_1585_),
    .X(_1586_));
 sky130_fd_sc_hd__o211ai_2 _6086_ (.A1(_1584_),
    .A2(_1585_),
    .B1(net154),
    .C1(_1424_),
    .Y(_1587_));
 sky130_fd_sc_hd__nand3_2 _6087_ (.A(_1480_),
    .B(_1586_),
    .C(_1587_),
    .Y(_1588_));
 sky130_fd_sc_hd__a21o_1 _6088_ (.A1(_1586_),
    .A2(_1587_),
    .B1(_1480_),
    .X(_1589_));
 sky130_fd_sc_hd__nand2_2 _6089_ (.A(_1588_),
    .B(_1589_),
    .Y(_1590_));
 sky130_fd_sc_hd__o21ba_2 _6090_ (.A1(_1323_),
    .A2(_1427_),
    .B1_N(_1426_),
    .X(_1591_));
 sky130_fd_sc_hd__xor2_4 _6091_ (.A(_1590_),
    .B(_1591_),
    .X(_1593_));
 sky130_fd_sc_hd__xnor2_4 _6092_ (.A(_1473_),
    .B(_1593_),
    .Y(_1594_));
 sky130_fd_sc_hd__and2b_1 _6093_ (.A_N(_1431_),
    .B(_1432_),
    .X(_1595_));
 sky130_fd_sc_hd__a21oi_4 _6094_ (.A1(_1319_),
    .A2(_1433_),
    .B1(_1595_),
    .Y(_1596_));
 sky130_fd_sc_hd__xnor2_4 _6095_ (.A(_1594_),
    .B(_1596_),
    .Y(_1597_));
 sky130_fd_sc_hd__or2_1 _6096_ (.A(_1435_),
    .B(_1434_),
    .X(_1598_));
 sky130_fd_sc_hd__and2_1 _6097_ (.A(_1597_),
    .B(_1598_),
    .X(_1599_));
 sky130_fd_sc_hd__nor2_1 _6098_ (.A(_1597_),
    .B(_1598_),
    .Y(_1600_));
 sky130_fd_sc_hd__or3_1 _6099_ (.A(_1138_),
    .B(_1265_),
    .C(_1434_),
    .X(_1601_));
 sky130_fd_sc_hd__o211ai_1 _6100_ (.A1(_1599_),
    .A2(_1600_),
    .B1(_1444_),
    .C1(_1601_),
    .Y(_1602_));
 sky130_fd_sc_hd__a211o_1 _6101_ (.A1(_1444_),
    .A2(_1601_),
    .B1(_1599_),
    .C1(_1600_),
    .X(_1604_));
 sky130_fd_sc_hd__and3_1 _6102_ (.A(_0320_),
    .B(_1602_),
    .C(_1604_),
    .X(_1605_));
 sky130_fd_sc_hd__a211o_1 _6103_ (.A1(_1458_),
    .A2(_1459_),
    .B1(_1472_),
    .C1(_1605_),
    .X(_1606_));
 sky130_fd_sc_hd__a31o_1 _6104_ (.A1(_3571_),
    .A2(_1453_),
    .A3(_1455_),
    .B1(_1606_),
    .X(net84));
 sky130_fd_sc_hd__buf_2 _6105_ (.A(net49),
    .X(_1607_));
 sky130_fd_sc_hd__clkbuf_4 _6106_ (.A(_1607_),
    .X(_1608_));
 sky130_fd_sc_hd__nor2_1 _6107_ (.A(_1756_),
    .B(_1608_),
    .Y(_1609_));
 sky130_fd_sc_hd__and2_1 _6108_ (.A(_1756_),
    .B(_1608_),
    .X(_1610_));
 sky130_fd_sc_hd__nor2_1 _6109_ (.A(_1609_),
    .B(_1610_),
    .Y(_1611_));
 sky130_fd_sc_hd__a21bo_1 _6110_ (.A1(_1297_),
    .A2(_1450_),
    .B1_N(_1451_),
    .X(_1612_));
 sky130_fd_sc_hd__a31o_1 _6111_ (.A1(_1456_),
    .A2(_1305_),
    .A3(_1452_),
    .B1(_1612_),
    .X(_1614_));
 sky130_fd_sc_hd__nand2_1 _6112_ (.A(_1611_),
    .B(_1614_),
    .Y(_1615_));
 sky130_fd_sc_hd__or2_1 _6113_ (.A(_1611_),
    .B(_1614_),
    .X(_1616_));
 sky130_fd_sc_hd__and3_1 _6114_ (.A(_0419_),
    .B(_1615_),
    .C(_1616_),
    .X(_1617_));
 sky130_fd_sc_hd__or3_1 _6115_ (.A(_1437_),
    .B(_1441_),
    .C(_1597_),
    .X(_1618_));
 sky130_fd_sc_hd__a311o_2 _6116_ (.A1(_0549_),
    .A2(_0552_),
    .A3(_0553_),
    .B1(_1145_),
    .C1(_1618_),
    .X(_1619_));
 sky130_fd_sc_hd__or2_2 _6117_ (.A(_1149_),
    .B(_1618_),
    .X(_1620_));
 sky130_fd_sc_hd__or2_1 _6118_ (.A(_1597_),
    .B(_1598_),
    .X(_1621_));
 sky130_fd_sc_hd__or3_1 _6119_ (.A(_1437_),
    .B(_1440_),
    .C(_1597_),
    .X(_1622_));
 sky130_fd_sc_hd__o211a_2 _6120_ (.A1(_1601_),
    .A2(_1599_),
    .B1(_1621_),
    .C1(_1622_),
    .X(_1623_));
 sky130_fd_sc_hd__and3_1 _6121_ (.A(net153),
    .B(_1620_),
    .C(_1623_),
    .X(_1625_));
 sky130_fd_sc_hd__or2_1 _6122_ (.A(_1594_),
    .B(_1596_),
    .X(_1626_));
 sky130_fd_sc_hd__or2_1 _6123_ (.A(_1590_),
    .B(_1591_),
    .X(_1627_));
 sky130_fd_sc_hd__a21bo_2 _6124_ (.A1(_1473_),
    .A2(_1593_),
    .B1_N(_1627_),
    .X(_1628_));
 sky130_fd_sc_hd__or2b_1 _6125_ (.A(_1495_),
    .B_N(_1496_),
    .X(_1629_));
 sky130_fd_sc_hd__or2_1 _6126_ (.A(_1488_),
    .B(_1497_),
    .X(_1630_));
 sky130_fd_sc_hd__o211a_1 _6127_ (.A1(_1483_),
    .A2(_1485_),
    .B1(_1384_),
    .C1(_1608_),
    .X(_1631_));
 sky130_fd_sc_hd__a211oi_1 _6128_ (.A1(_1384_),
    .A2(_1608_),
    .B1(_1483_),
    .C1(_1485_),
    .Y(_1632_));
 sky130_fd_sc_hd__or2_1 _6129_ (.A(_1631_),
    .B(_1632_),
    .X(_1633_));
 sky130_fd_sc_hd__a21oi_1 _6130_ (.A1(_1629_),
    .A2(_1630_),
    .B1(_1633_),
    .Y(_1634_));
 sky130_fd_sc_hd__and3_1 _6131_ (.A(_1629_),
    .B(_1630_),
    .C(_1633_),
    .X(_1636_));
 sky130_fd_sc_hd__nor2_1 _6132_ (.A(_1634_),
    .B(_1636_),
    .Y(_1637_));
 sky130_fd_sc_hd__xnor2_1 _6133_ (.A(_1475_),
    .B(_1637_),
    .Y(_1638_));
 sky130_fd_sc_hd__a21oi_1 _6134_ (.A1(_1516_),
    .A2(_1518_),
    .B1(_1638_),
    .Y(_1639_));
 sky130_fd_sc_hd__and3_1 _6135_ (.A(_1516_),
    .B(_1518_),
    .C(_1638_),
    .X(_1640_));
 sky130_fd_sc_hd__nor2_1 _6136_ (.A(_1639_),
    .B(_1640_),
    .Y(_1641_));
 sky130_fd_sc_hd__o211a_1 _6137_ (.A1(_1418_),
    .A2(net109),
    .B1(_1579_),
    .C1(_1580_),
    .X(_1642_));
 sky130_fd_sc_hd__inv_2 _6138_ (.A(_1511_),
    .Y(_1643_));
 sky130_fd_sc_hd__and3_1 _6139_ (.A(_1498_),
    .B(_1511_),
    .C(_1512_),
    .X(_1644_));
 sky130_fd_sc_hd__nand4_1 _6140_ (.A(_0215_),
    .B(_0346_),
    .C(_1169_),
    .D(_1294_),
    .Y(_1645_));
 sky130_fd_sc_hd__a22o_1 _6141_ (.A1(_0215_),
    .A2(_1169_),
    .B1(_1294_),
    .B2(_0346_),
    .X(_1647_));
 sky130_fd_sc_hd__nand2_1 _6142_ (.A(_1645_),
    .B(_1647_),
    .Y(_1648_));
 sky130_fd_sc_hd__nand2_1 _6143_ (.A(_1056_),
    .B(net48),
    .Y(_1649_));
 sky130_fd_sc_hd__xnor2_2 _6144_ (.A(_1648_),
    .B(_1649_),
    .Y(_1650_));
 sky130_fd_sc_hd__and4_1 _6145_ (.A(_2313_),
    .B(_2379_),
    .C(_0720_),
    .D(_0873_),
    .X(_1651_));
 sky130_fd_sc_hd__a22oi_1 _6146_ (.A1(_2379_),
    .A2(_0720_),
    .B1(_0873_),
    .B2(_2313_),
    .Y(_1652_));
 sky130_fd_sc_hd__and4bb_1 _6147_ (.A_N(_1651_),
    .B_N(_1652_),
    .C(_0106_),
    .D(net45),
    .X(_1653_));
 sky130_fd_sc_hd__o2bb2a_1 _6148_ (.A1_N(_0106_),
    .A2_N(_1007_),
    .B1(_1651_),
    .B2(_1652_),
    .X(_1654_));
 sky130_fd_sc_hd__nor2_1 _6149_ (.A(_1653_),
    .B(_1654_),
    .Y(_1655_));
 sky130_fd_sc_hd__or2_1 _6150_ (.A(_1489_),
    .B(_1491_),
    .X(_1656_));
 sky130_fd_sc_hd__xnor2_1 _6151_ (.A(_1655_),
    .B(_1656_),
    .Y(_1658_));
 sky130_fd_sc_hd__xor2_2 _6152_ (.A(_1650_),
    .B(_1658_),
    .X(_1659_));
 sky130_fd_sc_hd__nand2_1 _6153_ (.A(_1502_),
    .B(_1505_),
    .Y(_1660_));
 sky130_fd_sc_hd__a32o_1 _6154_ (.A1(_2160_),
    .A2(_0219_),
    .A3(_1524_),
    .B1(_1523_),
    .B2(_3719_),
    .X(_1661_));
 sky130_fd_sc_hd__nand4_1 _6155_ (.A(_2117_),
    .B(_2160_),
    .C(_0326_),
    .D(_0453_),
    .Y(_1662_));
 sky130_fd_sc_hd__a22o_1 _6156_ (.A1(_0247_),
    .A2(_0326_),
    .B1(_0453_),
    .B2(_2117_),
    .X(_1663_));
 sky130_fd_sc_hd__nand4_1 _6157_ (.A(_2445_),
    .B(_0688_),
    .C(_1662_),
    .D(_1663_),
    .Y(_1664_));
 sky130_fd_sc_hd__a22o_1 _6158_ (.A1(_2445_),
    .A2(_0688_),
    .B1(_1662_),
    .B2(_1663_),
    .X(_1665_));
 sky130_fd_sc_hd__nand3_1 _6159_ (.A(_1661_),
    .B(_1664_),
    .C(_1665_),
    .Y(_1666_));
 sky130_fd_sc_hd__a21o_1 _6160_ (.A1(_1664_),
    .A2(_1665_),
    .B1(_1661_),
    .X(_1667_));
 sky130_fd_sc_hd__nand3_1 _6161_ (.A(_1660_),
    .B(_1666_),
    .C(_1667_),
    .Y(_1669_));
 sky130_fd_sc_hd__a21o_1 _6162_ (.A1(_1666_),
    .A2(_1667_),
    .B1(_1660_),
    .X(_1670_));
 sky130_fd_sc_hd__a21o_1 _6163_ (.A1(_1500_),
    .A2(_1508_),
    .B1(_1507_),
    .X(_1671_));
 sky130_fd_sc_hd__nand3_1 _6164_ (.A(_1669_),
    .B(_1670_),
    .C(_1671_),
    .Y(_1672_));
 sky130_fd_sc_hd__a21o_1 _6165_ (.A1(_1669_),
    .A2(_1670_),
    .B1(_1671_),
    .X(_1673_));
 sky130_fd_sc_hd__nand3_2 _6166_ (.A(_1659_),
    .B(_1672_),
    .C(_1673_),
    .Y(_1674_));
 sky130_fd_sc_hd__a21o_1 _6167_ (.A1(_1672_),
    .A2(_1673_),
    .B1(_1659_),
    .X(_1675_));
 sky130_fd_sc_hd__o211ai_4 _6168_ (.A1(_1539_),
    .A2(_1541_),
    .B1(_1674_),
    .C1(_1675_),
    .Y(_1676_));
 sky130_fd_sc_hd__a211o_1 _6169_ (.A1(_1674_),
    .A2(_1675_),
    .B1(_1539_),
    .C1(_1541_),
    .X(_1677_));
 sky130_fd_sc_hd__o211a_1 _6170_ (.A1(_1643_),
    .A2(_1644_),
    .B1(_1676_),
    .C1(_1677_),
    .X(_1678_));
 sky130_fd_sc_hd__a211oi_2 _6171_ (.A1(_1676_),
    .A2(_1677_),
    .B1(_1643_),
    .C1(_1644_),
    .Y(_1680_));
 sky130_fd_sc_hd__a21o_1 _6172_ (.A1(_1544_),
    .A2(_1552_),
    .B1(_1551_),
    .X(_1681_));
 sky130_fd_sc_hd__a22o_1 _6173_ (.A1(_0491_),
    .A2(_0339_),
    .B1(_0099_),
    .B2(_2248_),
    .X(_1682_));
 sky130_fd_sc_hd__nand4_4 _6174_ (.A(_2248_),
    .B(_2653_),
    .C(_0339_),
    .D(_0099_),
    .Y(_1683_));
 sky130_fd_sc_hd__nand4_2 _6175_ (.A(_2215_),
    .B(_0219_),
    .C(_1682_),
    .D(_1683_),
    .Y(_1684_));
 sky130_fd_sc_hd__a22o_1 _6176_ (.A1(_2215_),
    .A2(_0219_),
    .B1(_1682_),
    .B2(_1683_),
    .X(_1685_));
 sky130_fd_sc_hd__and2_1 _6177_ (.A(_1684_),
    .B(_1685_),
    .X(_1686_));
 sky130_fd_sc_hd__nand4_2 _6178_ (.A(_0104_),
    .B(_3511_),
    .C(_2740_),
    .D(_0380_),
    .Y(_1687_));
 sky130_fd_sc_hd__a22o_1 _6179_ (.A1(_3511_),
    .A2(_2740_),
    .B1(_0380_),
    .B2(_3422_),
    .X(_1688_));
 sky130_fd_sc_hd__and4_2 _6180_ (.A(_3619_),
    .B(_2696_),
    .C(_1687_),
    .D(_1688_),
    .X(_1689_));
 sky130_fd_sc_hd__a22oi_4 _6181_ (.A1(_3620_),
    .A2(_2707_),
    .B1(_1687_),
    .B2(_1688_),
    .Y(_1691_));
 sky130_fd_sc_hd__a211o_2 _6182_ (.A1(_1530_),
    .A2(_1532_),
    .B1(_1689_),
    .C1(_1691_),
    .X(_1692_));
 sky130_fd_sc_hd__o211ai_4 _6183_ (.A1(_1689_),
    .A2(_1691_),
    .B1(_1530_),
    .C1(_1532_),
    .Y(_1693_));
 sky130_fd_sc_hd__nand3_4 _6184_ (.A(_1686_),
    .B(_1692_),
    .C(_1693_),
    .Y(_1694_));
 sky130_fd_sc_hd__a21o_1 _6185_ (.A1(_1692_),
    .A2(_1693_),
    .B1(_1686_),
    .X(_1695_));
 sky130_fd_sc_hd__and3_2 _6186_ (.A(_1681_),
    .B(_1694_),
    .C(_1695_),
    .X(_1696_));
 sky130_fd_sc_hd__a21oi_2 _6187_ (.A1(_1694_),
    .A2(_1695_),
    .B1(_1681_),
    .Y(_1697_));
 sky130_fd_sc_hd__a211oi_4 _6188_ (.A1(_1534_),
    .A2(_1536_),
    .B1(_1696_),
    .C1(_1697_),
    .Y(_1698_));
 sky130_fd_sc_hd__o211a_1 _6189_ (.A1(_1696_),
    .A2(_1697_),
    .B1(_1534_),
    .C1(_1536_),
    .X(_1699_));
 sky130_fd_sc_hd__nor3_1 _6190_ (.A(_1554_),
    .B(_1573_),
    .C(_1574_),
    .Y(_1700_));
 sky130_fd_sc_hd__nand4_2 _6191_ (.A(_0488_),
    .B(_0390_),
    .C(net16),
    .D(net17),
    .Y(_1702_));
 sky130_fd_sc_hd__a22o_1 _6192_ (.A1(net178),
    .A2(net16),
    .B1(net17),
    .B2(_3242_),
    .X(_1703_));
 sky130_fd_sc_hd__and2_1 _6193_ (.A(_0281_),
    .B(net15),
    .X(_1704_));
 sky130_fd_sc_hd__nand3_1 _6194_ (.A(_1702_),
    .B(_1703_),
    .C(_1704_),
    .Y(_1705_));
 sky130_fd_sc_hd__a21o_1 _6195_ (.A1(_1702_),
    .A2(_1703_),
    .B1(_1704_),
    .X(_1706_));
 sky130_fd_sc_hd__a21bo_1 _6196_ (.A1(_1556_),
    .A2(_1557_),
    .B1_N(_1555_),
    .X(_1707_));
 sky130_fd_sc_hd__nand3_1 _6197_ (.A(_1705_),
    .B(_1706_),
    .C(_1707_),
    .Y(_1708_));
 sky130_fd_sc_hd__a21o_1 _6198_ (.A1(_1705_),
    .A2(_1706_),
    .B1(_1707_),
    .X(_1709_));
 sky130_fd_sc_hd__and3_1 _6199_ (.A(_3169_),
    .B(net191),
    .C(net13),
    .X(_1710_));
 sky130_fd_sc_hd__a22o_1 _6200_ (.A1(_0030_),
    .A2(net13),
    .B1(net14),
    .B2(_3169_),
    .X(_1711_));
 sky130_fd_sc_hd__a21bo_1 _6201_ (.A1(_1887_),
    .A2(_1710_),
    .B1_N(_1711_),
    .X(_1713_));
 sky130_fd_sc_hd__nand2_1 _6202_ (.A(_2881_),
    .B(_2598_),
    .Y(_1714_));
 sky130_fd_sc_hd__xor2_1 _6203_ (.A(_1713_),
    .B(_1714_),
    .X(_1715_));
 sky130_fd_sc_hd__nand3_1 _6204_ (.A(_1708_),
    .B(_1709_),
    .C(_1715_),
    .Y(_1716_));
 sky130_fd_sc_hd__a21o_1 _6205_ (.A1(_1708_),
    .A2(_1709_),
    .B1(_1715_),
    .X(_1717_));
 sky130_fd_sc_hd__a21bo_1 _6206_ (.A1(_1563_),
    .A2(_1568_),
    .B1_N(_1562_),
    .X(_1718_));
 sky130_fd_sc_hd__and3_1 _6207_ (.A(_1716_),
    .B(_1717_),
    .C(_1718_),
    .X(_1719_));
 sky130_fd_sc_hd__clkbuf_2 _6208_ (.A(_1719_),
    .X(_1720_));
 sky130_fd_sc_hd__a21oi_2 _6209_ (.A1(_1716_),
    .A2(_1717_),
    .B1(_1718_),
    .Y(_1721_));
 sky130_fd_sc_hd__nand2_1 _6210_ (.A(_1546_),
    .B(_1549_),
    .Y(_1722_));
 sky130_fd_sc_hd__a32o_2 _6211_ (.A1(_2892_),
    .A2(_2576_),
    .A3(_1565_),
    .B1(_1564_),
    .B2(_1865_),
    .X(_1724_));
 sky130_fd_sc_hd__and4_1 _6212_ (.A(_3195_),
    .B(_3431_),
    .C(net9),
    .D(net10),
    .X(_1725_));
 sky130_fd_sc_hd__a22oi_2 _6213_ (.A1(_3271_),
    .A2(_2521_),
    .B1(_2565_),
    .B2(_3632_),
    .Y(_1726_));
 sky130_fd_sc_hd__and4bb_1 _6214_ (.A_N(_1725_),
    .B_N(_1726_),
    .C(_3430_),
    .D(_2499_),
    .X(_1727_));
 sky130_fd_sc_hd__o2bb2a_1 _6215_ (.A1_N(_3430_),
    .A2_N(_2499_),
    .B1(_1725_),
    .B2(_1726_),
    .X(_1728_));
 sky130_fd_sc_hd__or2_1 _6216_ (.A(_1727_),
    .B(_1728_),
    .X(_1729_));
 sky130_fd_sc_hd__xnor2_1 _6217_ (.A(_1724_),
    .B(_1729_),
    .Y(_1730_));
 sky130_fd_sc_hd__xnor2_1 _6218_ (.A(_1722_),
    .B(_1730_),
    .Y(_1731_));
 sky130_fd_sc_hd__or3_1 _6219_ (.A(_1720_),
    .B(_1721_),
    .C(_1731_),
    .X(_1732_));
 sky130_fd_sc_hd__o21ai_1 _6220_ (.A1(_1720_),
    .A2(_1721_),
    .B1(_1731_),
    .Y(_1733_));
 sky130_fd_sc_hd__o211a_2 _6221_ (.A1(_1573_),
    .A2(_1700_),
    .B1(_1732_),
    .C1(_1733_),
    .X(_1735_));
 sky130_fd_sc_hd__a211oi_1 _6222_ (.A1(_1732_),
    .A2(_1733_),
    .B1(_1573_),
    .C1(_1700_),
    .Y(_1736_));
 sky130_fd_sc_hd__nor4_1 _6223_ (.A(_1698_),
    .B(_1699_),
    .C(_1735_),
    .D(_1736_),
    .Y(_1737_));
 sky130_fd_sc_hd__o22a_1 _6224_ (.A1(_1698_),
    .A2(_1699_),
    .B1(_1735_),
    .B2(_1736_),
    .X(_1738_));
 sky130_fd_sc_hd__a211oi_4 _6225_ (.A1(_1577_),
    .A2(_1579_),
    .B1(net108),
    .C1(_1738_),
    .Y(_1739_));
 sky130_fd_sc_hd__o211a_1 _6226_ (.A1(net108),
    .A2(_1738_),
    .B1(_1577_),
    .C1(_1579_),
    .X(_1740_));
 sky130_fd_sc_hd__or4_1 _6227_ (.A(_1678_),
    .B(_1680_),
    .C(_1739_),
    .D(_1740_),
    .X(_1741_));
 sky130_fd_sc_hd__o22ai_2 _6228_ (.A1(_1678_),
    .A2(_1680_),
    .B1(_1739_),
    .B2(_1740_),
    .Y(_1742_));
 sky130_fd_sc_hd__o211ai_2 _6229_ (.A1(_1642_),
    .A2(_1584_),
    .B1(_1741_),
    .C1(_1742_),
    .Y(_1743_));
 sky130_fd_sc_hd__a211o_1 _6230_ (.A1(_1741_),
    .A2(_1742_),
    .B1(_1642_),
    .C1(_1584_),
    .X(_1744_));
 sky130_fd_sc_hd__and3_2 _6231_ (.A(_1641_),
    .B(_1743_),
    .C(_1744_),
    .X(_1746_));
 sky130_fd_sc_hd__a21oi_1 _6232_ (.A1(_1743_),
    .A2(_1744_),
    .B1(_1641_),
    .Y(_1747_));
 sky130_fd_sc_hd__a211oi_2 _6233_ (.A1(_1586_),
    .A2(_1588_),
    .B1(_1746_),
    .C1(_1747_),
    .Y(_1748_));
 sky130_fd_sc_hd__o211a_1 _6234_ (.A1(_1746_),
    .A2(_1747_),
    .B1(_1586_),
    .C1(_1588_),
    .X(_1749_));
 sky130_fd_sc_hd__nor3_1 _6235_ (.A(_1478_),
    .B(_1748_),
    .C(_1749_),
    .Y(_1750_));
 sky130_fd_sc_hd__o21a_1 _6236_ (.A1(_1748_),
    .A2(_1749_),
    .B1(_1478_),
    .X(_1751_));
 sky130_fd_sc_hd__nor2_2 _6237_ (.A(_1750_),
    .B(_1751_),
    .Y(_1752_));
 sky130_fd_sc_hd__xor2_4 _6238_ (.A(_1628_),
    .B(_1752_),
    .X(_1753_));
 sky130_fd_sc_hd__xor2_2 _6239_ (.A(_1626_),
    .B(_1753_),
    .X(_1754_));
 sky130_fd_sc_hd__o21a_1 _6240_ (.A1(_1625_),
    .A2(_1754_),
    .B1(_3305_),
    .X(_1755_));
 sky130_fd_sc_hd__a21boi_1 _6241_ (.A1(_1625_),
    .A2(_1754_),
    .B1_N(_1755_),
    .Y(_1757_));
 sky130_fd_sc_hd__mux4_1 _6242_ (.A0(_1756_),
    .A1(_1963_),
    .A2(_1942_),
    .A3(_1909_),
    .S0(_0583_),
    .S1(_0584_),
    .X(_1758_));
 sky130_fd_sc_hd__mux4_1 _6243_ (.A0(_0004_),
    .A1(_0585_),
    .A2(_1017_),
    .A3(_1758_),
    .S0(_0429_),
    .S1(_0189_),
    .X(_1759_));
 sky130_fd_sc_hd__nand2_1 _6244_ (.A(_0428_),
    .B(_3410_),
    .Y(_1760_));
 sky130_fd_sc_hd__o211a_1 _6245_ (.A1(_0428_),
    .A2(_1759_),
    .B1(_1760_),
    .C1(_0849_),
    .X(_1761_));
 sky130_fd_sc_hd__nor2_1 _6246_ (.A(_3156_),
    .B(_3404_),
    .Y(_1762_));
 sky130_fd_sc_hd__nand2_1 _6247_ (.A(_1756_),
    .B(_1608_),
    .Y(_1763_));
 sky130_fd_sc_hd__a21oi_1 _6248_ (.A1(_0438_),
    .A2(_1763_),
    .B1(_0000_),
    .Y(_1764_));
 sky130_fd_sc_hd__nor2_1 _6249_ (.A(_1609_),
    .B(_1764_),
    .Y(_1765_));
 sky130_fd_sc_hd__o31a_1 _6250_ (.A1(_0199_),
    .A2(_3727_),
    .A3(_3487_),
    .B1(_3161_),
    .X(_1766_));
 sky130_fd_sc_hd__a221o_1 _6251_ (.A1(_3414_),
    .A2(_1609_),
    .B1(_1610_),
    .B2(_0854_),
    .C1(_1766_),
    .X(_1768_));
 sky130_fd_sc_hd__or4_1 _6252_ (.A(_1761_),
    .B(_1762_),
    .C(_1765_),
    .D(_1768_),
    .X(_1769_));
 sky130_fd_sc_hd__or2_1 _6253_ (.A(_1609_),
    .B(_1610_),
    .X(_1770_));
 sky130_fd_sc_hd__and4_1 _6254_ (.A(_1011_),
    .B(_1272_),
    .C(_1299_),
    .D(_1454_),
    .X(_1771_));
 sky130_fd_sc_hd__and4_1 _6255_ (.A(_0563_),
    .B(_0693_),
    .C(_0829_),
    .D(_0878_),
    .X(_1772_));
 sky130_fd_sc_hd__inv_2 _6256_ (.A(_1448_),
    .Y(_1773_));
 sky130_fd_sc_hd__a21o_1 _6257_ (.A1(_0693_),
    .A2(_0694_),
    .B1(_0830_),
    .X(_1774_));
 sky130_fd_sc_hd__a21o_1 _6258_ (.A1(_0829_),
    .A2(_1774_),
    .B1(_1000_),
    .X(_1775_));
 sky130_fd_sc_hd__a21o_1 _6259_ (.A1(_0878_),
    .A2(_1775_),
    .B1(_1013_),
    .X(_1776_));
 sky130_fd_sc_hd__a21o_1 _6260_ (.A1(_1272_),
    .A2(_1273_),
    .B1(_1300_),
    .X(_1777_));
 sky130_fd_sc_hd__a21oi_1 _6261_ (.A1(_1299_),
    .A2(_1777_),
    .B1(_1446_),
    .Y(_1779_));
 sky130_fd_sc_hd__nor2_1 _6262_ (.A(_1452_),
    .B(_1779_),
    .Y(_1780_));
 sky130_fd_sc_hd__a221o_1 _6263_ (.A1(_1963_),
    .A2(_1773_),
    .B1(_1771_),
    .B2(_1776_),
    .C1(_1780_),
    .X(_1781_));
 sky130_fd_sc_hd__a31o_1 _6264_ (.A1(_0567_),
    .A2(_1771_),
    .A3(_1772_),
    .B1(_1781_),
    .X(_1782_));
 sky130_fd_sc_hd__a21oi_1 _6265_ (.A1(_1770_),
    .A2(_1782_),
    .B1(_0181_),
    .Y(_1783_));
 sky130_fd_sc_hd__o21a_1 _6266_ (.A1(_1770_),
    .A2(_1782_),
    .B1(_1783_),
    .X(_1784_));
 sky130_fd_sc_hd__or4_1 _6267_ (.A(_1617_),
    .B(_1757_),
    .C(_1769_),
    .D(_1784_),
    .X(_1785_));
 sky130_fd_sc_hd__buf_6 _6268_ (.A(_1785_),
    .X(net85));
 sky130_fd_sc_hd__or2b_1 _6269_ (.A(_1626_),
    .B_N(_1753_),
    .X(_1786_));
 sky130_fd_sc_hd__o21ai_1 _6270_ (.A1(_1625_),
    .A2(_1754_),
    .B1(_1786_),
    .Y(_1787_));
 sky130_fd_sc_hd__nand2_2 _6271_ (.A(_1628_),
    .B(_1752_),
    .Y(_1789_));
 sky130_fd_sc_hd__inv_2 _6272_ (.A(_1743_),
    .Y(_1790_));
 sky130_fd_sc_hd__nand2_1 _6273_ (.A(_1475_),
    .B(_1637_),
    .Y(_1791_));
 sky130_fd_sc_hd__o211ai_2 _6274_ (.A1(_1643_),
    .A2(_1644_),
    .B1(_1676_),
    .C1(_1677_),
    .Y(_1792_));
 sky130_fd_sc_hd__nand2_1 _6275_ (.A(_1676_),
    .B(_1792_),
    .Y(_1793_));
 sky130_fd_sc_hd__nand2_1 _6276_ (.A(_1655_),
    .B(_1656_),
    .Y(_1794_));
 sky130_fd_sc_hd__or2_1 _6277_ (.A(_1650_),
    .B(_1658_),
    .X(_1795_));
 sky130_fd_sc_hd__o21ai_1 _6278_ (.A1(_1648_),
    .A2(_1649_),
    .B1(_1645_),
    .Y(_1796_));
 sky130_fd_sc_hd__clkbuf_4 _6279_ (.A(net50),
    .X(_1797_));
 sky130_fd_sc_hd__a22oi_1 _6280_ (.A1(_1056_),
    .A2(_1607_),
    .B1(_1797_),
    .B2(_0991_),
    .Y(_1798_));
 sky130_fd_sc_hd__and4_1 _6281_ (.A(_0445_),
    .B(_0991_),
    .C(_1607_),
    .D(net50),
    .X(_1800_));
 sky130_fd_sc_hd__nor2_1 _6282_ (.A(_1798_),
    .B(_1800_),
    .Y(_1801_));
 sky130_fd_sc_hd__nand2_1 _6283_ (.A(_1796_),
    .B(_1801_),
    .Y(_1802_));
 sky130_fd_sc_hd__or2_1 _6284_ (.A(_1796_),
    .B(_1801_),
    .X(_1803_));
 sky130_fd_sc_hd__nand2_1 _6285_ (.A(_1802_),
    .B(_1803_),
    .Y(_1804_));
 sky130_fd_sc_hd__nand3_2 _6286_ (.A(_1794_),
    .B(_1795_),
    .C(_1804_),
    .Y(_1805_));
 sky130_fd_sc_hd__inv_2 _6287_ (.A(_1805_),
    .Y(_1806_));
 sky130_fd_sc_hd__a21oi_1 _6288_ (.A1(_1794_),
    .A2(_1795_),
    .B1(_1804_),
    .Y(_1807_));
 sky130_fd_sc_hd__or2_1 _6289_ (.A(_1806_),
    .B(_1807_),
    .X(_1808_));
 sky130_fd_sc_hd__nor2_1 _6290_ (.A(_1631_),
    .B(_1634_),
    .Y(_1809_));
 sky130_fd_sc_hd__xnor2_2 _6291_ (.A(_1808_),
    .B(_1809_),
    .Y(_1811_));
 sky130_fd_sc_hd__xnor2_1 _6292_ (.A(_1793_),
    .B(_1811_),
    .Y(_1812_));
 sky130_fd_sc_hd__xnor2_1 _6293_ (.A(_1791_),
    .B(_1812_),
    .Y(_1813_));
 sky130_fd_sc_hd__nor4_1 _6294_ (.A(_1678_),
    .B(_1680_),
    .C(_1739_),
    .D(_1740_),
    .Y(_1814_));
 sky130_fd_sc_hd__and2_1 _6295_ (.A(_1672_),
    .B(_1674_),
    .X(_1815_));
 sky130_fd_sc_hd__and4_1 _6296_ (.A(_0095_),
    .B(_0205_),
    .C(net46),
    .D(net47),
    .X(_1816_));
 sky130_fd_sc_hd__a22o_1 _6297_ (.A1(_0106_),
    .A2(net46),
    .B1(net47),
    .B2(_0205_),
    .X(_1817_));
 sky130_fd_sc_hd__or2b_1 _6298_ (.A(_1816_),
    .B_N(_1817_),
    .X(_1818_));
 sky130_fd_sc_hd__nand2_1 _6299_ (.A(_0357_),
    .B(net48),
    .Y(_1819_));
 sky130_fd_sc_hd__xnor2_1 _6300_ (.A(_1818_),
    .B(_1819_),
    .Y(_1820_));
 sky130_fd_sc_hd__nand4_2 _6301_ (.A(_2379_),
    .B(_2445_),
    .C(_0720_),
    .D(_0873_),
    .Y(_1822_));
 sky130_fd_sc_hd__a22o_1 _6302_ (.A1(_3530_),
    .A2(_0720_),
    .B1(_0873_),
    .B2(_2379_),
    .X(_1823_));
 sky130_fd_sc_hd__nand4_2 _6303_ (.A(_2324_),
    .B(_1007_),
    .C(_1822_),
    .D(_1823_),
    .Y(_1824_));
 sky130_fd_sc_hd__a22o_1 _6304_ (.A1(_2324_),
    .A2(net45),
    .B1(_1822_),
    .B2(_1823_),
    .X(_1825_));
 sky130_fd_sc_hd__o211ai_1 _6305_ (.A1(_1651_),
    .A2(_1653_),
    .B1(_1824_),
    .C1(_1825_),
    .Y(_1826_));
 sky130_fd_sc_hd__a211o_1 _6306_ (.A1(_1824_),
    .A2(_1825_),
    .B1(_1651_),
    .C1(_1653_),
    .X(_1827_));
 sky130_fd_sc_hd__nand2_1 _6307_ (.A(_1826_),
    .B(_1827_),
    .Y(_1828_));
 sky130_fd_sc_hd__xor2_1 _6308_ (.A(_1820_),
    .B(_1828_),
    .X(_1829_));
 sky130_fd_sc_hd__nand2_1 _6309_ (.A(_1662_),
    .B(_1664_),
    .Y(_1830_));
 sky130_fd_sc_hd__and4_1 _6310_ (.A(_0247_),
    .B(_2204_),
    .C(_0326_),
    .D(_0453_),
    .X(_1831_));
 sky130_fd_sc_hd__a22oi_1 _6311_ (.A1(_2204_),
    .A2(_0326_),
    .B1(_0453_),
    .B2(_0247_),
    .Y(_1833_));
 sky130_fd_sc_hd__and4bb_1 _6312_ (.A_N(_1831_),
    .B_N(_1833_),
    .C(_2117_),
    .D(_0654_),
    .X(_1834_));
 sky130_fd_sc_hd__o2bb2a_1 _6313_ (.A1_N(_2117_),
    .A2_N(_0654_),
    .B1(_1831_),
    .B2(_1833_),
    .X(_1835_));
 sky130_fd_sc_hd__a211o_1 _6314_ (.A1(_1683_),
    .A2(_1684_),
    .B1(_1834_),
    .C1(_1835_),
    .X(_1836_));
 sky130_fd_sc_hd__o211ai_2 _6315_ (.A1(_1834_),
    .A2(_1835_),
    .B1(_1683_),
    .C1(_1684_),
    .Y(_1837_));
 sky130_fd_sc_hd__nand3_2 _6316_ (.A(_1830_),
    .B(_1836_),
    .C(_1837_),
    .Y(_1838_));
 sky130_fd_sc_hd__a21o_1 _6317_ (.A1(_1836_),
    .A2(_1837_),
    .B1(_1830_),
    .X(_1839_));
 sky130_fd_sc_hd__a21bo_1 _6318_ (.A1(_1660_),
    .A2(_1667_),
    .B1_N(_1666_),
    .X(_1840_));
 sky130_fd_sc_hd__nand3_1 _6319_ (.A(_1838_),
    .B(_1839_),
    .C(_1840_),
    .Y(_1841_));
 sky130_fd_sc_hd__a21o_1 _6320_ (.A1(_1838_),
    .A2(_1839_),
    .B1(_1840_),
    .X(_1842_));
 sky130_fd_sc_hd__nand3_1 _6321_ (.A(_1829_),
    .B(_1841_),
    .C(_1842_),
    .Y(_1844_));
 sky130_fd_sc_hd__a21o_1 _6322_ (.A1(_1841_),
    .A2(_1842_),
    .B1(_1829_),
    .X(_1845_));
 sky130_fd_sc_hd__o211a_1 _6323_ (.A1(_1696_),
    .A2(_1698_),
    .B1(_1844_),
    .C1(_1845_),
    .X(_1846_));
 sky130_fd_sc_hd__a211o_1 _6324_ (.A1(_1844_),
    .A2(_1845_),
    .B1(_1696_),
    .C1(_1698_),
    .X(_1847_));
 sky130_fd_sc_hd__nor3b_2 _6325_ (.A(_1815_),
    .B(_1846_),
    .C_N(_1847_),
    .Y(_1848_));
 sky130_fd_sc_hd__or2b_1 _6326_ (.A(_1846_),
    .B_N(_1847_),
    .X(_1849_));
 sky130_fd_sc_hd__and2_1 _6327_ (.A(_1815_),
    .B(_1849_),
    .X(_1850_));
 sky130_fd_sc_hd__nor3_2 _6328_ (.A(_1720_),
    .B(_1721_),
    .C(_1731_),
    .Y(_1851_));
 sky130_fd_sc_hd__nand4_2 _6329_ (.A(_3451_),
    .B(_3452_),
    .C(net17),
    .D(net18),
    .Y(_1852_));
 sky130_fd_sc_hd__a22o_1 _6330_ (.A1(_0390_),
    .A2(net17),
    .B1(net18),
    .B2(_0488_),
    .X(_1853_));
 sky130_fd_sc_hd__and2_1 _6331_ (.A(_0292_),
    .B(net16),
    .X(_1855_));
 sky130_fd_sc_hd__nand3_1 _6332_ (.A(_1852_),
    .B(_1853_),
    .C(_1855_),
    .Y(_1856_));
 sky130_fd_sc_hd__a21o_1 _6333_ (.A1(_1852_),
    .A2(_1853_),
    .B1(_1855_),
    .X(_1857_));
 sky130_fd_sc_hd__a21bo_1 _6334_ (.A1(_1703_),
    .A2(_1704_),
    .B1_N(_1702_),
    .X(_1858_));
 sky130_fd_sc_hd__nand3_1 _6335_ (.A(_1856_),
    .B(_1857_),
    .C(_1858_),
    .Y(_1859_));
 sky130_fd_sc_hd__a21o_1 _6336_ (.A1(_1856_),
    .A2(_1857_),
    .B1(_1858_),
    .X(_1860_));
 sky130_fd_sc_hd__and3_1 _6337_ (.A(_3352_),
    .B(_0373_),
    .C(_1887_),
    .X(_1861_));
 sky130_fd_sc_hd__a22o_1 _6338_ (.A1(_0373_),
    .A2(_1887_),
    .B1(net15),
    .B2(_3352_),
    .X(_1862_));
 sky130_fd_sc_hd__a21bo_1 _6339_ (.A1(_1931_),
    .A2(_1861_),
    .B1_N(_1862_),
    .X(_1863_));
 sky130_fd_sc_hd__nand2_1 _6340_ (.A(_0042_),
    .B(_1854_),
    .Y(_1864_));
 sky130_fd_sc_hd__xor2_1 _6341_ (.A(_1863_),
    .B(_1864_),
    .X(_1866_));
 sky130_fd_sc_hd__nand3_1 _6342_ (.A(_1859_),
    .B(_1860_),
    .C(_1866_),
    .Y(_1867_));
 sky130_fd_sc_hd__a21o_1 _6343_ (.A1(_1859_),
    .A2(_1860_),
    .B1(_1866_),
    .X(_1868_));
 sky130_fd_sc_hd__a21bo_1 _6344_ (.A1(_1709_),
    .A2(_1715_),
    .B1_N(_1708_),
    .X(_1869_));
 sky130_fd_sc_hd__and3_2 _6345_ (.A(_1867_),
    .B(_1868_),
    .C(_1869_),
    .X(_1870_));
 sky130_fd_sc_hd__a21oi_2 _6346_ (.A1(_1867_),
    .A2(_1868_),
    .B1(_1869_),
    .Y(_1871_));
 sky130_fd_sc_hd__or2_1 _6347_ (.A(_1725_),
    .B(_1727_),
    .X(_1872_));
 sky130_fd_sc_hd__a32o_1 _6348_ (.A1(_2892_),
    .A2(_2598_),
    .A3(_1711_),
    .B1(_1710_),
    .B2(_1898_),
    .X(_1873_));
 sky130_fd_sc_hd__and4_1 _6349_ (.A(_3433_),
    .B(net162),
    .C(net10),
    .D(net11),
    .X(_1874_));
 sky130_fd_sc_hd__a22oi_1 _6350_ (.A1(_3633_),
    .A2(net10),
    .B1(net11),
    .B2(_3195_),
    .Y(_1875_));
 sky130_fd_sc_hd__and4bb_1 _6351_ (.A_N(_1874_),
    .B_N(_1875_),
    .C(_3343_),
    .D(_2521_),
    .X(_1877_));
 sky130_fd_sc_hd__o2bb2a_1 _6352_ (.A1_N(_3430_),
    .A2_N(_2532_),
    .B1(_1874_),
    .B2(_1875_),
    .X(_1878_));
 sky130_fd_sc_hd__or2_1 _6353_ (.A(_1877_),
    .B(_1878_),
    .X(_1879_));
 sky130_fd_sc_hd__xnor2_1 _6354_ (.A(_1873_),
    .B(_1879_),
    .Y(_1880_));
 sky130_fd_sc_hd__xnor2_1 _6355_ (.A(_1872_),
    .B(_1880_),
    .Y(_1881_));
 sky130_fd_sc_hd__or3_2 _6356_ (.A(_1870_),
    .B(_1871_),
    .C(_1881_),
    .X(_1882_));
 sky130_fd_sc_hd__o21ai_2 _6357_ (.A1(_1870_),
    .A2(_1871_),
    .B1(_1881_),
    .Y(_1883_));
 sky130_fd_sc_hd__o211a_1 _6358_ (.A1(_1720_),
    .A2(_1851_),
    .B1(_1882_),
    .C1(_1883_),
    .X(_1884_));
 sky130_fd_sc_hd__a211oi_2 _6359_ (.A1(_1882_),
    .A2(_1883_),
    .B1(_1720_),
    .C1(_1851_),
    .Y(_1885_));
 sky130_fd_sc_hd__and2b_1 _6360_ (.A_N(_1729_),
    .B(_1724_),
    .X(_1886_));
 sky130_fd_sc_hd__and2_1 _6361_ (.A(_1722_),
    .B(_1730_),
    .X(_1888_));
 sky130_fd_sc_hd__nand3_1 _6362_ (.A(_2707_),
    .B(_0100_),
    .C(_3722_),
    .Y(_1889_));
 sky130_fd_sc_hd__a22o_1 _6363_ (.A1(_3718_),
    .A2(_2696_),
    .B1(_0100_),
    .B2(_2653_),
    .X(_1890_));
 sky130_fd_sc_hd__nand4_1 _6364_ (.A(_2259_),
    .B(_0220_),
    .C(_1889_),
    .D(_1890_),
    .Y(_1891_));
 sky130_fd_sc_hd__a22o_1 _6365_ (.A1(_2259_),
    .A2(_0220_),
    .B1(_1889_),
    .B2(_1890_),
    .X(_1892_));
 sky130_fd_sc_hd__nand2_1 _6366_ (.A(_1891_),
    .B(_1892_),
    .Y(_1893_));
 sky130_fd_sc_hd__nand4_1 _6367_ (.A(_3423_),
    .B(_0105_),
    .C(_2773_),
    .D(_2499_),
    .Y(_1894_));
 sky130_fd_sc_hd__a22o_1 _6368_ (.A1(_0105_),
    .A2(_2773_),
    .B1(_2489_),
    .B2(_0104_),
    .X(_1895_));
 sky130_fd_sc_hd__nand2_1 _6369_ (.A(_1894_),
    .B(_1895_),
    .Y(_1896_));
 sky130_fd_sc_hd__and2_1 _6370_ (.A(_3619_),
    .B(_2751_),
    .X(_1897_));
 sky130_fd_sc_hd__xor2_1 _6371_ (.A(_1896_),
    .B(_1897_),
    .X(_1899_));
 sky130_fd_sc_hd__a41o_1 _6372_ (.A1(_3424_),
    .A2(_3512_),
    .A3(_2751_),
    .A4(_2773_),
    .B1(_1689_),
    .X(_1900_));
 sky130_fd_sc_hd__xor2_1 _6373_ (.A(_1899_),
    .B(_1900_),
    .X(_1901_));
 sky130_fd_sc_hd__xor2_1 _6374_ (.A(_1893_),
    .B(_1901_),
    .X(_1902_));
 sky130_fd_sc_hd__o21a_2 _6375_ (.A1(_1886_),
    .A2(_1888_),
    .B1(_1902_),
    .X(_1903_));
 sky130_fd_sc_hd__nor3_1 _6376_ (.A(_1886_),
    .B(_1888_),
    .C(_1902_),
    .Y(_1904_));
 sky130_fd_sc_hd__a211oi_4 _6377_ (.A1(_1692_),
    .A2(_1694_),
    .B1(_1903_),
    .C1(net120),
    .Y(_1905_));
 sky130_fd_sc_hd__o211a_1 _6378_ (.A1(_1903_),
    .A2(_1904_),
    .B1(_1692_),
    .C1(_1694_),
    .X(_1906_));
 sky130_fd_sc_hd__or4_4 _6379_ (.A(_1884_),
    .B(_1885_),
    .C(_1905_),
    .D(_1906_),
    .X(_1907_));
 sky130_fd_sc_hd__o22ai_4 _6380_ (.A1(_1884_),
    .A2(_1885_),
    .B1(_1905_),
    .B2(_1906_),
    .Y(_1908_));
 sky130_fd_sc_hd__o211a_2 _6381_ (.A1(_1735_),
    .A2(net201),
    .B1(_1907_),
    .C1(_1908_),
    .X(_1910_));
 sky130_fd_sc_hd__a211oi_4 _6382_ (.A1(_1907_),
    .A2(_1908_),
    .B1(_1735_),
    .C1(net201),
    .Y(_1911_));
 sky130_fd_sc_hd__or4_2 _6383_ (.A(_1848_),
    .B(_1850_),
    .C(_1910_),
    .D(_1911_),
    .X(_1912_));
 sky130_fd_sc_hd__o22ai_4 _6384_ (.A1(_1848_),
    .A2(_1850_),
    .B1(_1910_),
    .B2(_1911_),
    .Y(_1913_));
 sky130_fd_sc_hd__o211ai_4 _6385_ (.A1(_1739_),
    .A2(net105),
    .B1(_1912_),
    .C1(_1913_),
    .Y(_1914_));
 sky130_fd_sc_hd__a211o_1 _6386_ (.A1(_1912_),
    .A2(_1913_),
    .B1(_1739_),
    .C1(_1814_),
    .X(_1915_));
 sky130_fd_sc_hd__nand3_2 _6387_ (.A(_1813_),
    .B(_1914_),
    .C(net185),
    .Y(_1916_));
 sky130_fd_sc_hd__a21o_1 _6388_ (.A1(_1914_),
    .A2(_1915_),
    .B1(_1813_),
    .X(_1917_));
 sky130_fd_sc_hd__o211ai_2 _6389_ (.A1(_1790_),
    .A2(_1746_),
    .B1(_1916_),
    .C1(_1917_),
    .Y(_1918_));
 sky130_fd_sc_hd__a211o_1 _6390_ (.A1(_1916_),
    .A2(_1917_),
    .B1(_1790_),
    .C1(_1746_),
    .X(_1919_));
 sky130_fd_sc_hd__and3_1 _6391_ (.A(_1639_),
    .B(_1918_),
    .C(_1919_),
    .X(_1921_));
 sky130_fd_sc_hd__a21oi_1 _6392_ (.A1(_1918_),
    .A2(_1919_),
    .B1(_1639_),
    .Y(_1922_));
 sky130_fd_sc_hd__or2_2 _6393_ (.A(_1921_),
    .B(_1922_),
    .X(_1923_));
 sky130_fd_sc_hd__nor2_2 _6394_ (.A(_1748_),
    .B(_1750_),
    .Y(_1924_));
 sky130_fd_sc_hd__xor2_2 _6395_ (.A(_1923_),
    .B(_1924_),
    .X(_1925_));
 sky130_fd_sc_hd__xor2_1 _6396_ (.A(_1789_),
    .B(_1925_),
    .X(_1926_));
 sky130_fd_sc_hd__xnor2_1 _6397_ (.A(_1787_),
    .B(_1926_),
    .Y(_1927_));
 sky130_fd_sc_hd__nor2_1 _6398_ (.A(_1778_),
    .B(_1797_),
    .Y(_1928_));
 sky130_fd_sc_hd__and2_1 _6399_ (.A(_1778_),
    .B(_1797_),
    .X(_1929_));
 sky130_fd_sc_hd__or2_2 _6400_ (.A(_1928_),
    .B(_1929_),
    .X(_1930_));
 sky130_fd_sc_hd__a21oi_1 _6401_ (.A1(_1763_),
    .A2(_1615_),
    .B1(_1930_),
    .Y(_1932_));
 sky130_fd_sc_hd__a31o_1 _6402_ (.A1(_1763_),
    .A2(_1615_),
    .A3(_1930_),
    .B1(_3596_),
    .X(_1933_));
 sky130_fd_sc_hd__nor2_1 _6403_ (.A(_1932_),
    .B(_1933_),
    .Y(_1934_));
 sky130_fd_sc_hd__and2b_1 _6404_ (.A_N(_1608_),
    .B(_1756_),
    .X(_1935_));
 sky130_fd_sc_hd__a21o_1 _6405_ (.A1(_1770_),
    .A2(_1782_),
    .B1(_1935_),
    .X(_1936_));
 sky130_fd_sc_hd__nand2_1 _6406_ (.A(_1930_),
    .B(_1936_),
    .Y(_1937_));
 sky130_fd_sc_hd__or2_1 _6407_ (.A(_1930_),
    .B(_1936_),
    .X(_1938_));
 sky130_fd_sc_hd__mux4_1 _6408_ (.A0(_1778_),
    .A1(_1756_),
    .A2(_1963_),
    .A3(_1942_),
    .S0(_0583_),
    .S1(_0584_),
    .X(_1939_));
 sky130_fd_sc_hd__mux4_1 _6409_ (.A0(_0187_),
    .A1(_0710_),
    .A2(_1283_),
    .A3(_1939_),
    .S0(_0429_),
    .S1(_0189_),
    .X(_1940_));
 sky130_fd_sc_hd__nand2_1 _6410_ (.A(_0848_),
    .B(_3503_),
    .Y(_1941_));
 sky130_fd_sc_hd__o211a_1 _6411_ (.A1(_0848_),
    .A2(_1940_),
    .B1(_1941_),
    .C1(_0849_),
    .X(_1943_));
 sky130_fd_sc_hd__a22o_1 _6412_ (.A1(_0855_),
    .A2(_1928_),
    .B1(_1929_),
    .B2(_0854_),
    .X(_1944_));
 sky130_fd_sc_hd__o21ba_1 _6413_ (.A1(_3589_),
    .A2(_1929_),
    .B1_N(_0000_),
    .X(_1945_));
 sky130_fd_sc_hd__o22a_1 _6414_ (.A1(_3156_),
    .A2(_3493_),
    .B1(_1928_),
    .B2(_1945_),
    .X(_1946_));
 sky130_fd_sc_hd__or4b_1 _6415_ (.A(_1766_),
    .B(_1943_),
    .C(_1944_),
    .D_N(_1946_),
    .X(_1947_));
 sky130_fd_sc_hd__a31o_1 _6416_ (.A1(_3571_),
    .A2(_1937_),
    .A3(_1938_),
    .B1(_1947_),
    .X(_1948_));
 sky130_fd_sc_hd__a211o_2 _6417_ (.A1(_0320_),
    .A2(_1927_),
    .B1(_1934_),
    .C1(_1948_),
    .X(net86));
 sky130_fd_sc_hd__buf_2 _6418_ (.A(net51),
    .X(_1949_));
 sky130_fd_sc_hd__nor2_1 _6419_ (.A(_1810_),
    .B(_1949_),
    .Y(_1950_));
 sky130_fd_sc_hd__and2_1 _6420_ (.A(_1810_),
    .B(_1949_),
    .X(_1951_));
 sky130_fd_sc_hd__or2_2 _6421_ (.A(_1950_),
    .B(_1951_),
    .X(_1953_));
 sky130_fd_sc_hd__o21bai_2 _6422_ (.A1(_1610_),
    .A2(_1929_),
    .B1_N(_1928_),
    .Y(_1954_));
 sky130_fd_sc_hd__nor2_1 _6423_ (.A(_1770_),
    .B(_1930_),
    .Y(_1955_));
 sky130_fd_sc_hd__nand2_1 _6424_ (.A(_1614_),
    .B(_1955_),
    .Y(_1956_));
 sky130_fd_sc_hd__nand3_1 _6425_ (.A(_1953_),
    .B(_1954_),
    .C(_1956_),
    .Y(_1957_));
 sky130_fd_sc_hd__a21o_1 _6426_ (.A1(_1954_),
    .A2(_1956_),
    .B1(_1953_),
    .X(_1958_));
 sky130_fd_sc_hd__and2b_1 _6427_ (.A_N(_1797_),
    .B(_1778_),
    .X(_1959_));
 sky130_fd_sc_hd__a21o_1 _6428_ (.A1(_1930_),
    .A2(_1936_),
    .B1(_1959_),
    .X(_1960_));
 sky130_fd_sc_hd__a21oi_1 _6429_ (.A1(_1953_),
    .A2(_1960_),
    .B1(_0181_),
    .Y(_1961_));
 sky130_fd_sc_hd__o21a_1 _6430_ (.A1(_1953_),
    .A2(_1960_),
    .B1(_1961_),
    .X(_1962_));
 sky130_fd_sc_hd__nor2_2 _6431_ (.A(_1923_),
    .B(_1924_),
    .Y(_1964_));
 sky130_fd_sc_hd__inv_2 _6432_ (.A(_1918_),
    .Y(_1965_));
 sky130_fd_sc_hd__a21oi_2 _6433_ (.A1(_1676_),
    .A2(_1792_),
    .B1(_1811_),
    .Y(_1966_));
 sky130_fd_sc_hd__and3_1 _6434_ (.A(_1475_),
    .B(_1637_),
    .C(_1812_),
    .X(_1967_));
 sky130_fd_sc_hd__or2_1 _6435_ (.A(_1846_),
    .B(_1848_),
    .X(_1968_));
 sky130_fd_sc_hd__o21ai_1 _6436_ (.A1(_1820_),
    .A2(_1828_),
    .B1(_1826_),
    .Y(_1969_));
 sky130_fd_sc_hd__a31o_1 _6437_ (.A1(_0357_),
    .A2(net48),
    .A3(_1817_),
    .B1(_1816_),
    .X(_1970_));
 sky130_fd_sc_hd__and4_1 _6438_ (.A(_0346_),
    .B(_0434_),
    .C(net49),
    .D(net50),
    .X(_1971_));
 sky130_fd_sc_hd__a22oi_1 _6439_ (.A1(_0346_),
    .A2(_1607_),
    .B1(net50),
    .B2(_0707_),
    .Y(_1972_));
 sky130_fd_sc_hd__and4bb_1 _6440_ (.A_N(_1971_),
    .B_N(_1972_),
    .C(_0991_),
    .D(net51),
    .X(_1973_));
 sky130_fd_sc_hd__o2bb2a_1 _6441_ (.A1_N(_0991_),
    .A2_N(net51),
    .B1(_1971_),
    .B2(_1972_),
    .X(_1975_));
 sky130_fd_sc_hd__or2_1 _6442_ (.A(_1973_),
    .B(_1975_),
    .X(_1976_));
 sky130_fd_sc_hd__xnor2_1 _6443_ (.A(_1970_),
    .B(_1976_),
    .Y(_1977_));
 sky130_fd_sc_hd__xnor2_1 _6444_ (.A(_1800_),
    .B(_1977_),
    .Y(_1978_));
 sky130_fd_sc_hd__xor2_1 _6445_ (.A(_1969_),
    .B(_1978_),
    .X(_1979_));
 sky130_fd_sc_hd__xor2_1 _6446_ (.A(_1802_),
    .B(_1979_),
    .X(_1980_));
 sky130_fd_sc_hd__or2_1 _6447_ (.A(_1631_),
    .B(_1807_),
    .X(_1981_));
 sky130_fd_sc_hd__nand3_2 _6448_ (.A(_1805_),
    .B(_1980_),
    .C(_1981_),
    .Y(_1982_));
 sky130_fd_sc_hd__a21o_1 _6449_ (.A1(_1805_),
    .A2(_1981_),
    .B1(_1980_),
    .X(_1983_));
 sky130_fd_sc_hd__and2_1 _6450_ (.A(_1982_),
    .B(_1983_),
    .X(_1984_));
 sky130_fd_sc_hd__xnor2_1 _6451_ (.A(_1968_),
    .B(_1984_),
    .Y(_1986_));
 sky130_fd_sc_hd__and3b_1 _6452_ (.A_N(_1807_),
    .B(_1634_),
    .C(_1805_),
    .X(_1987_));
 sky130_fd_sc_hd__xnor2_1 _6453_ (.A(_1986_),
    .B(_1987_),
    .Y(_1988_));
 sky130_fd_sc_hd__nor4_1 _6454_ (.A(_1848_),
    .B(_1850_),
    .C(_1910_),
    .D(_1911_),
    .Y(_1989_));
 sky130_fd_sc_hd__o211ai_2 _6455_ (.A1(_1720_),
    .A2(_1851_),
    .B1(_1882_),
    .C1(_1883_),
    .Y(_1990_));
 sky130_fd_sc_hd__nor3_1 _6456_ (.A(_1870_),
    .B(_1871_),
    .C(_1881_),
    .Y(_1991_));
 sky130_fd_sc_hd__nand4_1 _6457_ (.A(_0499_),
    .B(_0401_),
    .C(_1767_),
    .D(_1799_),
    .Y(_1992_));
 sky130_fd_sc_hd__a22o_1 _6458_ (.A1(_0401_),
    .A2(_1767_),
    .B1(net19),
    .B2(_0499_),
    .X(_1993_));
 sky130_fd_sc_hd__and2_1 _6459_ (.A(_0303_),
    .B(net17),
    .X(_1994_));
 sky130_fd_sc_hd__nand3_1 _6460_ (.A(_1992_),
    .B(_1993_),
    .C(_1994_),
    .Y(_1995_));
 sky130_fd_sc_hd__a21o_1 _6461_ (.A1(_1992_),
    .A2(_1993_),
    .B1(_1994_),
    .X(_1997_));
 sky130_fd_sc_hd__a21bo_1 _6462_ (.A1(_1853_),
    .A2(_1855_),
    .B1_N(_1852_),
    .X(_1998_));
 sky130_fd_sc_hd__nand3_1 _6463_ (.A(_1995_),
    .B(_1997_),
    .C(_1998_),
    .Y(_1999_));
 sky130_fd_sc_hd__a21o_1 _6464_ (.A1(_1995_),
    .A2(_1997_),
    .B1(_1998_),
    .X(_2000_));
 sky130_fd_sc_hd__and3_1 _6465_ (.A(_3645_),
    .B(_0041_),
    .C(net15),
    .X(_2001_));
 sky130_fd_sc_hd__a22o_1 _6466_ (.A1(_0041_),
    .A2(net15),
    .B1(net16),
    .B2(_3645_),
    .X(_2002_));
 sky130_fd_sc_hd__a21bo_1 _6467_ (.A1(_1952_),
    .A2(_2001_),
    .B1_N(_2002_),
    .X(_2003_));
 sky130_fd_sc_hd__nand2_1 _6468_ (.A(_2892_),
    .B(_1898_),
    .Y(_2004_));
 sky130_fd_sc_hd__xor2_1 _6469_ (.A(_2003_),
    .B(_2004_),
    .X(_2005_));
 sky130_fd_sc_hd__nand3_1 _6470_ (.A(_1999_),
    .B(_2000_),
    .C(_2005_),
    .Y(_2006_));
 sky130_fd_sc_hd__a21o_1 _6471_ (.A1(_1999_),
    .A2(_2000_),
    .B1(_2005_),
    .X(_2008_));
 sky130_fd_sc_hd__a21bo_1 _6472_ (.A1(_1860_),
    .A2(_1866_),
    .B1_N(_1859_),
    .X(_2009_));
 sky130_fd_sc_hd__and3_1 _6473_ (.A(_2006_),
    .B(_2008_),
    .C(_2009_),
    .X(_2010_));
 sky130_fd_sc_hd__buf_2 _6474_ (.A(_2010_),
    .X(_2011_));
 sky130_fd_sc_hd__a21oi_2 _6475_ (.A1(_2006_),
    .A2(_2008_),
    .B1(_2009_),
    .Y(_2012_));
 sky130_fd_sc_hd__or2_2 _6476_ (.A(_1874_),
    .B(_1877_),
    .X(_2013_));
 sky130_fd_sc_hd__a32o_1 _6477_ (.A1(_2892_),
    .A2(_1865_),
    .A3(_1862_),
    .B1(_1861_),
    .B2(_1931_),
    .X(_2014_));
 sky130_fd_sc_hd__and4_1 _6478_ (.A(_3196_),
    .B(_3272_),
    .C(_2598_),
    .D(_1854_),
    .X(_2015_));
 sky130_fd_sc_hd__a22oi_1 _6479_ (.A1(_3272_),
    .A2(_2598_),
    .B1(_1854_),
    .B2(_3196_),
    .Y(_2016_));
 sky130_fd_sc_hd__and4bb_1 _6480_ (.A_N(_2015_),
    .B_N(_2016_),
    .C(_3385_),
    .D(_2576_),
    .X(_2017_));
 sky130_fd_sc_hd__o2bb2a_1 _6481_ (.A1_N(_3385_),
    .A2_N(_2576_),
    .B1(_2015_),
    .B2(_2016_),
    .X(_2019_));
 sky130_fd_sc_hd__or2_1 _6482_ (.A(_2017_),
    .B(_2019_),
    .X(_2020_));
 sky130_fd_sc_hd__xnor2_2 _6483_ (.A(_2014_),
    .B(_2020_),
    .Y(_2021_));
 sky130_fd_sc_hd__xnor2_2 _6484_ (.A(_2013_),
    .B(_2021_),
    .Y(_2022_));
 sky130_fd_sc_hd__or3_2 _6485_ (.A(_2011_),
    .B(_2012_),
    .C(_2022_),
    .X(_2023_));
 sky130_fd_sc_hd__o21ai_2 _6486_ (.A1(_2011_),
    .A2(_2012_),
    .B1(_2022_),
    .Y(_2024_));
 sky130_fd_sc_hd__o211a_1 _6487_ (.A1(_1870_),
    .A2(_1991_),
    .B1(_2023_),
    .C1(_2024_),
    .X(_2025_));
 sky130_fd_sc_hd__a211oi_1 _6488_ (.A1(_2023_),
    .A2(_2024_),
    .B1(_1870_),
    .C1(_1991_),
    .Y(_2026_));
 sky130_fd_sc_hd__or2b_1 _6489_ (.A(_1899_),
    .B_N(_1900_),
    .X(_2027_));
 sky130_fd_sc_hd__or2_1 _6490_ (.A(_1893_),
    .B(_1901_),
    .X(_2028_));
 sky130_fd_sc_hd__and2b_1 _6491_ (.A_N(_1879_),
    .B(_1873_),
    .X(_2030_));
 sky130_fd_sc_hd__and2_1 _6492_ (.A(_1872_),
    .B(_1880_),
    .X(_2031_));
 sky130_fd_sc_hd__a21o_1 _6493_ (.A1(_3720_),
    .A2(_2751_),
    .B1(_0191_),
    .X(_2032_));
 sky130_fd_sc_hd__nand3_1 _6494_ (.A(_3720_),
    .B(_2762_),
    .C(_0191_),
    .Y(_2033_));
 sky130_fd_sc_hd__nand2_1 _6495_ (.A(_2032_),
    .B(_2033_),
    .Y(_2034_));
 sky130_fd_sc_hd__nor2_1 _6496_ (.A(_0178_),
    .B(_0337_),
    .Y(_2035_));
 sky130_fd_sc_hd__xor2_2 _6497_ (.A(_2034_),
    .B(_2035_),
    .X(_2036_));
 sky130_fd_sc_hd__nand4_1 _6498_ (.A(_3424_),
    .B(_3512_),
    .C(_2499_),
    .D(_2532_),
    .Y(_2037_));
 sky130_fd_sc_hd__a22o_1 _6499_ (.A1(_3512_),
    .A2(_2499_),
    .B1(_2532_),
    .B2(_3423_),
    .X(_2038_));
 sky130_fd_sc_hd__and4_1 _6500_ (.A(_3620_),
    .B(_2784_),
    .C(_2037_),
    .D(_2038_),
    .X(_2039_));
 sky130_fd_sc_hd__a22oi_1 _6501_ (.A1(_3620_),
    .A2(_2784_),
    .B1(_2037_),
    .B2(_2038_),
    .Y(_2041_));
 sky130_fd_sc_hd__a21bo_1 _6502_ (.A1(_1895_),
    .A2(_1897_),
    .B1_N(_1894_),
    .X(_2042_));
 sky130_fd_sc_hd__or3b_2 _6503_ (.A(_2039_),
    .B(_2041_),
    .C_N(_2042_),
    .X(_2043_));
 sky130_fd_sc_hd__o21bai_1 _6504_ (.A1(_2039_),
    .A2(_2041_),
    .B1_N(_2042_),
    .Y(_2044_));
 sky130_fd_sc_hd__nand2_1 _6505_ (.A(_2043_),
    .B(_2044_),
    .Y(_2045_));
 sky130_fd_sc_hd__xor2_2 _6506_ (.A(_2036_),
    .B(_2045_),
    .X(_2046_));
 sky130_fd_sc_hd__o21a_1 _6507_ (.A1(_2030_),
    .A2(_2031_),
    .B1(_2046_),
    .X(_2047_));
 sky130_fd_sc_hd__nor3_1 _6508_ (.A(_2030_),
    .B(_2031_),
    .C(_2046_),
    .Y(_2048_));
 sky130_fd_sc_hd__a211oi_2 _6509_ (.A1(_2027_),
    .A2(_2028_),
    .B1(_2047_),
    .C1(_2048_),
    .Y(_2049_));
 sky130_fd_sc_hd__o211a_1 _6510_ (.A1(_2047_),
    .A2(_2048_),
    .B1(_2027_),
    .C1(_2028_),
    .X(_2050_));
 sky130_fd_sc_hd__nor4_1 _6511_ (.A(_2025_),
    .B(_2026_),
    .C(_2049_),
    .D(_2050_),
    .Y(_2052_));
 sky130_fd_sc_hd__o22a_1 _6512_ (.A1(_2025_),
    .A2(_2026_),
    .B1(_2049_),
    .B2(_2050_),
    .X(_2053_));
 sky130_fd_sc_hd__a211oi_2 _6513_ (.A1(_1990_),
    .A2(_1907_),
    .B1(net200),
    .C1(_2053_),
    .Y(_2054_));
 sky130_fd_sc_hd__o211a_1 _6514_ (.A1(_2052_),
    .A2(_2053_),
    .B1(_1990_),
    .C1(_1907_),
    .X(_2055_));
 sky130_fd_sc_hd__nand2_1 _6515_ (.A(_1841_),
    .B(_1844_),
    .Y(_2056_));
 sky130_fd_sc_hd__nand4_2 _6516_ (.A(_0117_),
    .B(_2335_),
    .C(_1170_),
    .D(_1295_),
    .Y(_2057_));
 sky130_fd_sc_hd__a22o_1 _6517_ (.A1(_2324_),
    .A2(_1169_),
    .B1(_1295_),
    .B2(_0106_),
    .X(_2058_));
 sky130_fd_sc_hd__nand4_1 _6518_ (.A(_0226_),
    .B(net48),
    .C(_2057_),
    .D(_2058_),
    .Y(_2059_));
 sky130_fd_sc_hd__a22o_1 _6519_ (.A1(_1034_),
    .A2(_1448_),
    .B1(_2057_),
    .B2(_2058_),
    .X(_2060_));
 sky130_fd_sc_hd__nand2_2 _6520_ (.A(_2059_),
    .B(_2060_),
    .Y(_2061_));
 sky130_fd_sc_hd__and4_1 _6521_ (.A(_2445_),
    .B(_2127_),
    .C(_0721_),
    .D(_0874_),
    .X(_2063_));
 sky130_fd_sc_hd__a22o_1 _6522_ (.A1(_2127_),
    .A2(_0721_),
    .B1(_0874_),
    .B2(_2445_),
    .X(_2064_));
 sky130_fd_sc_hd__or2b_1 _6523_ (.A(_2063_),
    .B_N(_2064_),
    .X(_2065_));
 sky130_fd_sc_hd__nand2_1 _6524_ (.A(_2401_),
    .B(_1007_),
    .Y(_2066_));
 sky130_fd_sc_hd__xnor2_2 _6525_ (.A(_2065_),
    .B(_2066_),
    .Y(_2067_));
 sky130_fd_sc_hd__nand2_1 _6526_ (.A(_1822_),
    .B(_1824_),
    .Y(_2068_));
 sky130_fd_sc_hd__xor2_2 _6527_ (.A(_2067_),
    .B(_2068_),
    .X(_2069_));
 sky130_fd_sc_hd__xor2_2 _6528_ (.A(_2061_),
    .B(_2069_),
    .X(_2070_));
 sky130_fd_sc_hd__or2_1 _6529_ (.A(_1831_),
    .B(_1834_),
    .X(_2071_));
 sky130_fd_sc_hd__and3_1 _6530_ (.A(_2707_),
    .B(_0100_),
    .C(_3722_),
    .X(_2072_));
 sky130_fd_sc_hd__a31o_1 _6531_ (.A1(_2270_),
    .A2(_0293_),
    .A3(_1890_),
    .B1(_2072_),
    .X(_2074_));
 sky130_fd_sc_hd__and4_1 _6532_ (.A(_2215_),
    .B(_2259_),
    .C(_0327_),
    .D(_0454_),
    .X(_2075_));
 sky130_fd_sc_hd__a22oi_1 _6533_ (.A1(_2259_),
    .A2(_0327_),
    .B1(_0454_),
    .B2(_2226_),
    .Y(_2076_));
 sky130_fd_sc_hd__and4bb_1 _6534_ (.A_N(_2075_),
    .B_N(_2076_),
    .C(_2160_),
    .D(_0688_),
    .X(_2077_));
 sky130_fd_sc_hd__o2bb2a_1 _6535_ (.A1_N(_2160_),
    .A2_N(_0688_),
    .B1(_2075_),
    .B2(_2076_),
    .X(_2078_));
 sky130_fd_sc_hd__or2_1 _6536_ (.A(_2077_),
    .B(_2078_),
    .X(_2079_));
 sky130_fd_sc_hd__xnor2_2 _6537_ (.A(_2074_),
    .B(_2079_),
    .Y(_2080_));
 sky130_fd_sc_hd__xnor2_1 _6538_ (.A(_2071_),
    .B(_2080_),
    .Y(_2081_));
 sky130_fd_sc_hd__a21o_1 _6539_ (.A1(_1836_),
    .A2(_1838_),
    .B1(_2081_),
    .X(_2082_));
 sky130_fd_sc_hd__nand3_1 _6540_ (.A(_1836_),
    .B(_1838_),
    .C(_2081_),
    .Y(_2083_));
 sky130_fd_sc_hd__nand3_2 _6541_ (.A(_2070_),
    .B(_2082_),
    .C(_2083_),
    .Y(_2085_));
 sky130_fd_sc_hd__a21o_1 _6542_ (.A1(_2082_),
    .A2(_2083_),
    .B1(_2070_),
    .X(_2086_));
 sky130_fd_sc_hd__o211ai_2 _6543_ (.A1(_1903_),
    .A2(_1905_),
    .B1(_2085_),
    .C1(_2086_),
    .Y(_2087_));
 sky130_fd_sc_hd__a211o_1 _6544_ (.A1(_2085_),
    .A2(_2086_),
    .B1(_1903_),
    .C1(_1905_),
    .X(_2088_));
 sky130_fd_sc_hd__nand3_1 _6545_ (.A(_2056_),
    .B(_2087_),
    .C(_2088_),
    .Y(_2089_));
 sky130_fd_sc_hd__a21o_1 _6546_ (.A1(_2087_),
    .A2(_2088_),
    .B1(_2056_),
    .X(_2090_));
 sky130_fd_sc_hd__or4bb_2 _6547_ (.A(_2054_),
    .B(_2055_),
    .C_N(_2089_),
    .D_N(_2090_),
    .X(_2091_));
 sky130_fd_sc_hd__a2bb2o_1 _6548_ (.A1_N(_2054_),
    .A2_N(_2055_),
    .B1(_2089_),
    .B2(_2090_),
    .X(_2092_));
 sky130_fd_sc_hd__o211ai_4 _6549_ (.A1(_1910_),
    .A2(net103),
    .B1(_2091_),
    .C1(_2092_),
    .Y(_2093_));
 sky130_fd_sc_hd__a211o_1 _6550_ (.A1(_2091_),
    .A2(_2092_),
    .B1(_1910_),
    .C1(_1989_),
    .X(_2094_));
 sky130_fd_sc_hd__and3_1 _6551_ (.A(_1988_),
    .B(_2093_),
    .C(_2094_),
    .X(_2096_));
 sky130_fd_sc_hd__a21oi_2 _6552_ (.A1(_2093_),
    .A2(net182),
    .B1(_1988_),
    .Y(_2097_));
 sky130_fd_sc_hd__a211o_1 _6553_ (.A1(_1914_),
    .A2(_1916_),
    .B1(_2096_),
    .C1(_2097_),
    .X(_2098_));
 sky130_fd_sc_hd__o211ai_4 _6554_ (.A1(net169),
    .A2(_2097_),
    .B1(_1914_),
    .C1(_1916_),
    .Y(_2099_));
 sky130_fd_sc_hd__o211ai_4 _6555_ (.A1(_1966_),
    .A2(_1967_),
    .B1(net157),
    .C1(_2099_),
    .Y(_2100_));
 sky130_fd_sc_hd__a211o_1 _6556_ (.A1(_2098_),
    .A2(_2099_),
    .B1(_1966_),
    .C1(_1967_),
    .X(_2101_));
 sky130_fd_sc_hd__o211ai_4 _6557_ (.A1(_1965_),
    .A2(net175),
    .B1(_2100_),
    .C1(net171),
    .Y(_2102_));
 sky130_fd_sc_hd__a211o_1 _6558_ (.A1(_2100_),
    .A2(_2101_),
    .B1(_1965_),
    .C1(net174),
    .X(_2103_));
 sky130_fd_sc_hd__and2_2 _6559_ (.A(_2102_),
    .B(_2103_),
    .X(_2104_));
 sky130_fd_sc_hd__xnor2_4 _6560_ (.A(_1964_),
    .B(_2104_),
    .Y(_2105_));
 sky130_fd_sc_hd__a21bo_1 _6561_ (.A1(_1789_),
    .A2(_1786_),
    .B1_N(_1925_),
    .X(_2107_));
 sky130_fd_sc_hd__or2_1 _6562_ (.A(_1754_),
    .B(_1926_),
    .X(_2108_));
 sky130_fd_sc_hd__a31o_1 _6563_ (.A1(_1619_),
    .A2(_1620_),
    .A3(_1623_),
    .B1(_2108_),
    .X(_2109_));
 sky130_fd_sc_hd__and3_1 _6564_ (.A(_2105_),
    .B(_2107_),
    .C(_2109_),
    .X(_2110_));
 sky130_fd_sc_hd__a21o_1 _6565_ (.A1(_2107_),
    .A2(_2109_),
    .B1(_2105_),
    .X(_2111_));
 sky130_fd_sc_hd__and3b_1 _6566_ (.A_N(_2110_),
    .B(_2111_),
    .C(_0320_),
    .X(_2112_));
 sky130_fd_sc_hd__a311o_1 _6567_ (.A1(_0419_),
    .A2(_1957_),
    .A3(_1958_),
    .B1(_1962_),
    .C1(_2112_),
    .X(_2113_));
 sky130_fd_sc_hd__mux4_1 _6568_ (.A0(_1810_),
    .A1(_1778_),
    .A2(_1756_),
    .A3(_1963_),
    .S0(_0863_),
    .S1(_0864_),
    .X(_2114_));
 sky130_fd_sc_hd__mux4_1 _6569_ (.A0(_0304_),
    .A1(_0845_),
    .A2(_1308_),
    .A3(_2114_),
    .S0(_0866_),
    .S1(_0867_),
    .X(_2115_));
 sky130_fd_sc_hd__nand2_1 _6570_ (.A(_0861_),
    .B(_3605_),
    .Y(_2116_));
 sky130_fd_sc_hd__o211a_1 _6571_ (.A1(_0861_),
    .A2(_2115_),
    .B1(_2116_),
    .C1(_0844_),
    .X(_2118_));
 sky130_fd_sc_hd__nand2_1 _6572_ (.A(_1810_),
    .B(_1949_),
    .Y(_2119_));
 sky130_fd_sc_hd__a21oi_1 _6573_ (.A1(_0438_),
    .A2(_2119_),
    .B1(_1277_),
    .Y(_2120_));
 sky130_fd_sc_hd__o31a_1 _6574_ (.A1(_0199_),
    .A2(_0428_),
    .A3(_3707_),
    .B1(_3161_),
    .X(_2121_));
 sky130_fd_sc_hd__a221o_1 _6575_ (.A1(_0855_),
    .A2(_1950_),
    .B1(_1951_),
    .B2(_0854_),
    .C1(_2121_),
    .X(_2122_));
 sky130_fd_sc_hd__o21ba_1 _6576_ (.A1(_1950_),
    .A2(_2120_),
    .B1_N(_2122_),
    .X(_2123_));
 sky130_fd_sc_hd__o21a_1 _6577_ (.A1(_3156_),
    .A2(_3585_),
    .B1(_2123_),
    .X(_2124_));
 sky130_fd_sc_hd__or3b_1 _6578_ (.A(_2113_),
    .B(_2118_),
    .C_N(_2124_),
    .X(_2125_));
 sky130_fd_sc_hd__clkbuf_2 _6579_ (.A(_2125_),
    .X(net87));
 sky130_fd_sc_hd__nand2_2 _6580_ (.A(_1964_),
    .B(_2104_),
    .Y(_2126_));
 sky130_fd_sc_hd__nand2_2 _6581_ (.A(net158),
    .B(_2100_),
    .Y(_2128_));
 sky130_fd_sc_hd__or2_1 _6582_ (.A(_1968_),
    .B(_1984_),
    .X(_2129_));
 sky130_fd_sc_hd__and2_1 _6583_ (.A(_1968_),
    .B(_1984_),
    .X(_2130_));
 sky130_fd_sc_hd__a21oi_2 _6584_ (.A1(_2129_),
    .A2(_1987_),
    .B1(_2130_),
    .Y(_2131_));
 sky130_fd_sc_hd__nor3_2 _6585_ (.A(_2011_),
    .B(_2012_),
    .C(_2022_),
    .Y(_2132_));
 sky130_fd_sc_hd__nand4_1 _6586_ (.A(_0499_),
    .B(_0401_),
    .C(_1799_),
    .D(net20),
    .Y(_2133_));
 sky130_fd_sc_hd__a22o_1 _6587_ (.A1(_0401_),
    .A2(_1799_),
    .B1(net20),
    .B2(_0499_),
    .X(_2134_));
 sky130_fd_sc_hd__and2_1 _6588_ (.A(_0303_),
    .B(_1767_),
    .X(_2135_));
 sky130_fd_sc_hd__nand3_1 _6589_ (.A(_2133_),
    .B(_2134_),
    .C(_2135_),
    .Y(_2136_));
 sky130_fd_sc_hd__a21o_1 _6590_ (.A1(_2133_),
    .A2(_2134_),
    .B1(_2135_),
    .X(_2137_));
 sky130_fd_sc_hd__a21bo_1 _6591_ (.A1(_1993_),
    .A2(_1994_),
    .B1_N(_1992_),
    .X(_2139_));
 sky130_fd_sc_hd__nand3_1 _6592_ (.A(_2136_),
    .B(_2137_),
    .C(_2139_),
    .Y(_2140_));
 sky130_fd_sc_hd__a21o_1 _6593_ (.A1(_2136_),
    .A2(_2137_),
    .B1(_2139_),
    .X(_2141_));
 sky130_fd_sc_hd__and3_1 _6594_ (.A(_0172_),
    .B(_0052_),
    .C(net16),
    .X(_2142_));
 sky130_fd_sc_hd__a22o_1 _6595_ (.A1(_0052_),
    .A2(net16),
    .B1(net17),
    .B2(_0172_),
    .X(_2143_));
 sky130_fd_sc_hd__a21bo_1 _6596_ (.A1(_1745_),
    .A2(_2142_),
    .B1_N(_2143_),
    .X(_2144_));
 sky130_fd_sc_hd__nand2_1 _6597_ (.A(_2892_),
    .B(_1931_),
    .Y(_2145_));
 sky130_fd_sc_hd__xor2_1 _6598_ (.A(_2144_),
    .B(_2145_),
    .X(_2146_));
 sky130_fd_sc_hd__nand3_1 _6599_ (.A(_2140_),
    .B(_2141_),
    .C(_2146_),
    .Y(_2147_));
 sky130_fd_sc_hd__a21o_1 _6600_ (.A1(_2140_),
    .A2(_2141_),
    .B1(_2146_),
    .X(_2148_));
 sky130_fd_sc_hd__a21bo_1 _6601_ (.A1(_2000_),
    .A2(_2005_),
    .B1_N(_1999_),
    .X(_2150_));
 sky130_fd_sc_hd__and3_2 _6602_ (.A(_2147_),
    .B(_2148_),
    .C(_2150_),
    .X(_2151_));
 sky130_fd_sc_hd__a21oi_2 _6603_ (.A1(net152),
    .A2(_2148_),
    .B1(_2150_),
    .Y(_2152_));
 sky130_fd_sc_hd__or2_1 _6604_ (.A(_2015_),
    .B(_2017_),
    .X(_2153_));
 sky130_fd_sc_hd__o2bb2a_1 _6605_ (.A1_N(_1952_),
    .A2_N(_2001_),
    .B1(_2003_),
    .B2(_2004_),
    .X(_2154_));
 sky130_fd_sc_hd__and4_1 _6606_ (.A(_3196_),
    .B(_3271_),
    .C(_1854_),
    .D(_1887_),
    .X(_2155_));
 sky130_fd_sc_hd__a22oi_1 _6607_ (.A1(_3272_),
    .A2(_1854_),
    .B1(_1898_),
    .B2(_3196_),
    .Y(_2156_));
 sky130_fd_sc_hd__and4bb_1 _6608_ (.A_N(_2155_),
    .B_N(_2156_),
    .C(_3385_),
    .D(_2598_),
    .X(_2157_));
 sky130_fd_sc_hd__o2bb2a_1 _6609_ (.A1_N(_3385_),
    .A2_N(_2609_),
    .B1(_2155_),
    .B2(_2156_),
    .X(_2158_));
 sky130_fd_sc_hd__or2_1 _6610_ (.A(_2157_),
    .B(_2158_),
    .X(_2159_));
 sky130_fd_sc_hd__xor2_2 _6611_ (.A(_2154_),
    .B(_2159_),
    .X(_2161_));
 sky130_fd_sc_hd__xnor2_2 _6612_ (.A(_2153_),
    .B(_2161_),
    .Y(_2162_));
 sky130_fd_sc_hd__or3_2 _6613_ (.A(_2151_),
    .B(_2152_),
    .C(_2162_),
    .X(_2163_));
 sky130_fd_sc_hd__o21ai_4 _6614_ (.A1(_2151_),
    .A2(_2152_),
    .B1(_2162_),
    .Y(_2164_));
 sky130_fd_sc_hd__o211a_1 _6615_ (.A1(_2011_),
    .A2(_2132_),
    .B1(_2163_),
    .C1(_2164_),
    .X(_2165_));
 sky130_fd_sc_hd__a211oi_2 _6616_ (.A1(_2163_),
    .A2(_2164_),
    .B1(_2011_),
    .C1(_2132_),
    .Y(_2166_));
 sky130_fd_sc_hd__or2_1 _6617_ (.A(_2036_),
    .B(_2045_),
    .X(_2167_));
 sky130_fd_sc_hd__and2b_1 _6618_ (.A_N(_2020_),
    .B(_2014_),
    .X(_2168_));
 sky130_fd_sc_hd__and2_1 _6619_ (.A(_2013_),
    .B(_2021_),
    .X(_2169_));
 sky130_fd_sc_hd__a22o_1 _6620_ (.A1(_0174_),
    .A2(_2751_),
    .B1(_2784_),
    .B2(_3719_),
    .X(_2170_));
 sky130_fd_sc_hd__nand4_2 _6621_ (.A(_3720_),
    .B(_0174_),
    .C(_2762_),
    .D(_2784_),
    .Y(_2172_));
 sky130_fd_sc_hd__a22o_1 _6622_ (.A1(_2718_),
    .A2(_0293_),
    .B1(_2170_),
    .B2(_2172_),
    .X(_2173_));
 sky130_fd_sc_hd__nand4_2 _6623_ (.A(_2718_),
    .B(_0293_),
    .C(_2170_),
    .D(_2172_),
    .Y(_2174_));
 sky130_fd_sc_hd__nand2_1 _6624_ (.A(_2173_),
    .B(_2174_),
    .Y(_2175_));
 sky130_fd_sc_hd__and4_1 _6625_ (.A(_3423_),
    .B(_3512_),
    .C(_2532_),
    .D(_2565_),
    .X(_2176_));
 sky130_fd_sc_hd__a22o_1 _6626_ (.A1(_3512_),
    .A2(_2532_),
    .B1(_2565_),
    .B2(_3423_),
    .X(_2177_));
 sky130_fd_sc_hd__or2b_1 _6627_ (.A(_2176_),
    .B_N(_2177_),
    .X(_2178_));
 sky130_fd_sc_hd__nand2_1 _6628_ (.A(_3620_),
    .B(_2510_),
    .Y(_2179_));
 sky130_fd_sc_hd__xnor2_1 _6629_ (.A(_2178_),
    .B(_2179_),
    .Y(_2180_));
 sky130_fd_sc_hd__a41o_1 _6630_ (.A1(_3425_),
    .A2(_3513_),
    .A3(_2510_),
    .A4(_2543_),
    .B1(_2039_),
    .X(_2181_));
 sky130_fd_sc_hd__xor2_1 _6631_ (.A(_2180_),
    .B(_2181_),
    .X(_2183_));
 sky130_fd_sc_hd__xor2_1 _6632_ (.A(_2175_),
    .B(_2183_),
    .X(_2184_));
 sky130_fd_sc_hd__o21a_2 _6633_ (.A1(_2168_),
    .A2(_2169_),
    .B1(_2184_),
    .X(_2185_));
 sky130_fd_sc_hd__nor3_1 _6634_ (.A(_2168_),
    .B(_2169_),
    .C(_2184_),
    .Y(_2186_));
 sky130_fd_sc_hd__a211oi_4 _6635_ (.A1(_2043_),
    .A2(_2167_),
    .B1(_2185_),
    .C1(net117),
    .Y(_2187_));
 sky130_fd_sc_hd__o211a_1 _6636_ (.A1(_2185_),
    .A2(_2186_),
    .B1(_2043_),
    .C1(_2167_),
    .X(_2188_));
 sky130_fd_sc_hd__or4_4 _6637_ (.A(_2165_),
    .B(_2166_),
    .C(_2187_),
    .D(_2188_),
    .X(_2189_));
 sky130_fd_sc_hd__o22ai_2 _6638_ (.A1(_2165_),
    .A2(_2166_),
    .B1(_2187_),
    .B2(_2188_),
    .Y(_2190_));
 sky130_fd_sc_hd__o211a_1 _6639_ (.A1(net189),
    .A2(net104),
    .B1(_2189_),
    .C1(_2190_),
    .X(_2191_));
 sky130_fd_sc_hd__a211oi_2 _6640_ (.A1(_2189_),
    .A2(_2190_),
    .B1(net189),
    .C1(net104),
    .Y(_2192_));
 sky130_fd_sc_hd__inv_2 _6641_ (.A(_2082_),
    .Y(_2194_));
 sky130_fd_sc_hd__and3_1 _6642_ (.A(_2070_),
    .B(_2082_),
    .C(_2083_),
    .X(_2195_));
 sky130_fd_sc_hd__inv_2 _6643_ (.A(net143),
    .Y(_2196_));
 sky130_fd_sc_hd__a211o_2 _6644_ (.A1(_2027_),
    .A2(_2028_),
    .B1(_2047_),
    .C1(_2048_),
    .X(_2197_));
 sky130_fd_sc_hd__a22o_1 _6645_ (.A1(_2390_),
    .A2(_1169_),
    .B1(_1294_),
    .B2(_2324_),
    .X(_2198_));
 sky130_fd_sc_hd__nand4_2 _6646_ (.A(_2324_),
    .B(_2390_),
    .C(_1169_),
    .D(_1294_),
    .Y(_2199_));
 sky130_fd_sc_hd__a22o_1 _6647_ (.A1(_0117_),
    .A2(net48),
    .B1(_2198_),
    .B2(_2199_),
    .X(_2200_));
 sky130_fd_sc_hd__nand4_2 _6648_ (.A(_0117_),
    .B(net48),
    .C(_2198_),
    .D(_2199_),
    .Y(_2201_));
 sky130_fd_sc_hd__nand2_1 _6649_ (.A(_2200_),
    .B(_2201_),
    .Y(_2202_));
 sky130_fd_sc_hd__nand4_1 _6650_ (.A(_2117_),
    .B(_2160_),
    .C(_0721_),
    .D(_0874_),
    .Y(_2203_));
 sky130_fd_sc_hd__a22o_1 _6651_ (.A1(_2160_),
    .A2(_0721_),
    .B1(_0874_),
    .B2(_2117_),
    .X(_2205_));
 sky130_fd_sc_hd__nand2_1 _6652_ (.A(_2203_),
    .B(_2205_),
    .Y(_2206_));
 sky130_fd_sc_hd__and2_1 _6653_ (.A(_2445_),
    .B(_1007_),
    .X(_2207_));
 sky130_fd_sc_hd__xor2_1 _6654_ (.A(_2206_),
    .B(_2207_),
    .X(_2208_));
 sky130_fd_sc_hd__a31o_1 _6655_ (.A1(_2401_),
    .A2(_1007_),
    .A3(_2064_),
    .B1(_2063_),
    .X(_2209_));
 sky130_fd_sc_hd__xor2_1 _6656_ (.A(_2208_),
    .B(_2209_),
    .X(_2210_));
 sky130_fd_sc_hd__or2_1 _6657_ (.A(_2202_),
    .B(_2210_),
    .X(_2211_));
 sky130_fd_sc_hd__nand2_1 _6658_ (.A(_2202_),
    .B(_2210_),
    .Y(_2212_));
 sky130_fd_sc_hd__and2_1 _6659_ (.A(_2211_),
    .B(_2212_),
    .X(_2213_));
 sky130_fd_sc_hd__or2b_1 _6660_ (.A(_2079_),
    .B_N(_2074_),
    .X(_2214_));
 sky130_fd_sc_hd__nand2_1 _6661_ (.A(_2071_),
    .B(_2080_),
    .Y(_2216_));
 sky130_fd_sc_hd__or2_1 _6662_ (.A(_2075_),
    .B(_2077_),
    .X(_2217_));
 sky130_fd_sc_hd__a21boi_2 _6663_ (.A1(_2032_),
    .A2(_2035_),
    .B1_N(_2033_),
    .Y(_2218_));
 sky130_fd_sc_hd__and4_1 _6664_ (.A(_2259_),
    .B(_2653_),
    .C(_0326_),
    .D(_0453_),
    .X(_2219_));
 sky130_fd_sc_hd__a22oi_1 _6665_ (.A1(_2664_),
    .A2(_0327_),
    .B1(_0454_),
    .B2(_2259_),
    .Y(_2220_));
 sky130_fd_sc_hd__and4bb_1 _6666_ (.A_N(_2219_),
    .B_N(_2220_),
    .C(_2226_),
    .D(_0688_),
    .X(_2221_));
 sky130_fd_sc_hd__o2bb2a_1 _6667_ (.A1_N(_2226_),
    .A2_N(_0688_),
    .B1(_2219_),
    .B2(_2220_),
    .X(_2222_));
 sky130_fd_sc_hd__or2_1 _6668_ (.A(_2221_),
    .B(_2222_),
    .X(_2223_));
 sky130_fd_sc_hd__xor2_2 _6669_ (.A(_2218_),
    .B(_2223_),
    .X(_2224_));
 sky130_fd_sc_hd__xnor2_2 _6670_ (.A(_2217_),
    .B(_2224_),
    .Y(_2225_));
 sky130_fd_sc_hd__a21o_1 _6671_ (.A1(_2214_),
    .A2(_2216_),
    .B1(_2225_),
    .X(_2227_));
 sky130_fd_sc_hd__nand3_1 _6672_ (.A(_2214_),
    .B(_2216_),
    .C(_2225_),
    .Y(_2228_));
 sky130_fd_sc_hd__and3_2 _6673_ (.A(_2213_),
    .B(_2227_),
    .C(_2228_),
    .X(_2229_));
 sky130_fd_sc_hd__a21oi_2 _6674_ (.A1(_2227_),
    .A2(_2228_),
    .B1(_2213_),
    .Y(_2230_));
 sky130_fd_sc_hd__a211o_2 _6675_ (.A1(_2196_),
    .A2(_2197_),
    .B1(_2229_),
    .C1(_2230_),
    .X(_2231_));
 sky130_fd_sc_hd__o211ai_4 _6676_ (.A1(_2229_),
    .A2(_2230_),
    .B1(_2196_),
    .C1(_2197_),
    .Y(_2232_));
 sky130_fd_sc_hd__o211ai_4 _6677_ (.A1(_2194_),
    .A2(_2195_),
    .B1(_2231_),
    .C1(_2232_),
    .Y(_2233_));
 sky130_fd_sc_hd__a211o_1 _6678_ (.A1(_2231_),
    .A2(_2232_),
    .B1(_2194_),
    .C1(_2195_),
    .X(_2234_));
 sky130_fd_sc_hd__and4bb_1 _6679_ (.A_N(_2191_),
    .B_N(_2192_),
    .C(_2233_),
    .D(_2234_),
    .X(_2235_));
 sky130_fd_sc_hd__a2bb2o_1 _6680_ (.A1_N(_2191_),
    .A2_N(_2192_),
    .B1(_2233_),
    .B2(_2234_),
    .X(_2236_));
 sky130_fd_sc_hd__or2b_1 _6681_ (.A(_2235_),
    .B_N(_2236_),
    .X(_2238_));
 sky130_fd_sc_hd__and2b_1 _6682_ (.A_N(_2054_),
    .B(_2091_),
    .X(_2239_));
 sky130_fd_sc_hd__xnor2_1 _6683_ (.A(_2238_),
    .B(_2239_),
    .Y(_2240_));
 sky130_fd_sc_hd__nand2_1 _6684_ (.A(_2087_),
    .B(_2089_),
    .Y(_2241_));
 sky130_fd_sc_hd__or2b_1 _6685_ (.A(_2067_),
    .B_N(_2068_),
    .X(_2242_));
 sky130_fd_sc_hd__o21ai_2 _6686_ (.A1(_2061_),
    .A2(_2069_),
    .B1(_2242_),
    .Y(_2243_));
 sky130_fd_sc_hd__or2_1 _6687_ (.A(_1971_),
    .B(_1973_),
    .X(_2244_));
 sky130_fd_sc_hd__nand2_1 _6688_ (.A(_2057_),
    .B(_2059_),
    .Y(_2245_));
 sky130_fd_sc_hd__a22o_1 _6689_ (.A1(_0205_),
    .A2(net49),
    .B1(net50),
    .B2(_0335_),
    .X(_2246_));
 sky130_fd_sc_hd__inv_2 _6690_ (.A(_2246_),
    .Y(_2247_));
 sky130_fd_sc_hd__and4_1 _6691_ (.A(_0215_),
    .B(_0346_),
    .C(_1607_),
    .D(net50),
    .X(_2249_));
 sky130_fd_sc_hd__o2bb2a_1 _6692_ (.A1_N(_1056_),
    .A2_N(net51),
    .B1(_2247_),
    .B2(_2249_),
    .X(_2250_));
 sky130_fd_sc_hd__and4b_1 _6693_ (.A_N(_2249_),
    .B(net51),
    .C(_1056_),
    .D(_2246_),
    .X(_2251_));
 sky130_fd_sc_hd__or2_1 _6694_ (.A(_2250_),
    .B(_2251_),
    .X(_2252_));
 sky130_fd_sc_hd__xnor2_1 _6695_ (.A(_2245_),
    .B(_2252_),
    .Y(_2253_));
 sky130_fd_sc_hd__xnor2_1 _6696_ (.A(_2244_),
    .B(_2253_),
    .Y(_2254_));
 sky130_fd_sc_hd__xor2_1 _6697_ (.A(_2243_),
    .B(_2254_),
    .X(_2255_));
 sky130_fd_sc_hd__and2b_1 _6698_ (.A_N(_1976_),
    .B(_1970_),
    .X(_2256_));
 sky130_fd_sc_hd__a21oi_1 _6699_ (.A1(_1800_),
    .A2(_1977_),
    .B1(_2256_),
    .Y(_2257_));
 sky130_fd_sc_hd__xnor2_1 _6700_ (.A(_2255_),
    .B(_2257_),
    .Y(_2258_));
 sky130_fd_sc_hd__and2b_1 _6701_ (.A_N(_1978_),
    .B(_1969_),
    .X(_2260_));
 sky130_fd_sc_hd__o21ba_1 _6702_ (.A1(_1802_),
    .A2(_1979_),
    .B1_N(_2260_),
    .X(_2261_));
 sky130_fd_sc_hd__xor2_1 _6703_ (.A(_2258_),
    .B(_2261_),
    .X(_2262_));
 sky130_fd_sc_hd__clkbuf_4 _6704_ (.A(net52),
    .X(_2263_));
 sky130_fd_sc_hd__nand2_1 _6705_ (.A(_3209_),
    .B(_2263_),
    .Y(_2264_));
 sky130_fd_sc_hd__xor2_1 _6706_ (.A(_2262_),
    .B(_2264_),
    .X(_2265_));
 sky130_fd_sc_hd__xnor2_1 _6707_ (.A(_2241_),
    .B(_2265_),
    .Y(_2266_));
 sky130_fd_sc_hd__xnor2_1 _6708_ (.A(_1982_),
    .B(_2266_),
    .Y(_2267_));
 sky130_fd_sc_hd__xnor2_1 _6709_ (.A(_2240_),
    .B(_2267_),
    .Y(_2268_));
 sky130_fd_sc_hd__inv_2 _6710_ (.A(_2093_),
    .Y(_2269_));
 sky130_fd_sc_hd__nor2_1 _6711_ (.A(_2269_),
    .B(net170),
    .Y(_2271_));
 sky130_fd_sc_hd__xnor2_1 _6712_ (.A(_2268_),
    .B(_2271_),
    .Y(_2272_));
 sky130_fd_sc_hd__xnor2_2 _6713_ (.A(_2131_),
    .B(_2272_),
    .Y(_2273_));
 sky130_fd_sc_hd__xnor2_4 _6714_ (.A(_2128_),
    .B(_2273_),
    .Y(_2274_));
 sky130_fd_sc_hd__xnor2_2 _6715_ (.A(_2102_),
    .B(_2274_),
    .Y(_2275_));
 sky130_fd_sc_hd__a21oi_1 _6716_ (.A1(_2126_),
    .A2(net177),
    .B1(_2275_),
    .Y(_2276_));
 sky130_fd_sc_hd__a311o_1 _6717_ (.A1(_2126_),
    .A2(net177),
    .A3(_2275_),
    .B1(_2276_),
    .C1(_3192_),
    .X(_2277_));
 sky130_fd_sc_hd__or2_2 _6718_ (.A(_1821_),
    .B(_2263_),
    .X(_2278_));
 sky130_fd_sc_hd__nand2_1 _6719_ (.A(_1821_),
    .B(_2263_),
    .Y(_2279_));
 sky130_fd_sc_hd__nand2_2 _6720_ (.A(_2278_),
    .B(_2279_),
    .Y(_2280_));
 sky130_fd_sc_hd__a21oi_1 _6721_ (.A1(_2119_),
    .A2(_1958_),
    .B1(_2280_),
    .Y(_2282_));
 sky130_fd_sc_hd__a31o_1 _6722_ (.A1(_2119_),
    .A2(_1958_),
    .A3(_2280_),
    .B1(_3596_),
    .X(_2283_));
 sky130_fd_sc_hd__or2_1 _6723_ (.A(_2282_),
    .B(_2283_),
    .X(_2284_));
 sky130_fd_sc_hd__mux4_1 _6724_ (.A0(_1821_),
    .A1(_1810_),
    .A2(_1778_),
    .A3(_1756_),
    .S0(_0863_),
    .S1(_0864_),
    .X(_2285_));
 sky130_fd_sc_hd__mux4_1 _6725_ (.A0(_0433_),
    .A1(_0865_),
    .A2(_1466_),
    .A3(_2285_),
    .S0(_0866_),
    .S1(_0867_),
    .X(_2286_));
 sky130_fd_sc_hd__nor2_1 _6726_ (.A(_0861_),
    .B(_2286_),
    .Y(_2287_));
 sky130_fd_sc_hd__a211o_1 _6727_ (.A1(_0861_),
    .A2(_3705_),
    .B1(_2287_),
    .C1(_3118_),
    .X(_2288_));
 sky130_fd_sc_hd__and2_1 _6728_ (.A(_0438_),
    .B(_2279_),
    .X(_2289_));
 sky130_fd_sc_hd__o21ai_1 _6729_ (.A1(_1277_),
    .A2(_2289_),
    .B1(_2278_),
    .Y(_2290_));
 sky130_fd_sc_hd__o22a_1 _6730_ (.A1(_3712_),
    .A2(_2278_),
    .B1(_2279_),
    .B2(_0309_),
    .X(_2291_));
 sky130_fd_sc_hd__and2b_1 _6731_ (.A_N(_2121_),
    .B(_2291_),
    .X(_2293_));
 sky130_fd_sc_hd__o2111a_1 _6732_ (.A1(_3156_),
    .A2(_3699_),
    .B1(_2288_),
    .C1(_2290_),
    .D1(_2293_),
    .X(_2294_));
 sky130_fd_sc_hd__and2b_1 _6733_ (.A_N(_1949_),
    .B(_1810_),
    .X(_2295_));
 sky130_fd_sc_hd__a21o_1 _6734_ (.A1(_1953_),
    .A2(_1960_),
    .B1(_2295_),
    .X(_2296_));
 sky130_fd_sc_hd__a21oi_1 _6735_ (.A1(_2280_),
    .A2(_2296_),
    .B1(_0181_),
    .Y(_2297_));
 sky130_fd_sc_hd__o21ai_1 _6736_ (.A1(_2280_),
    .A2(_2296_),
    .B1(_2297_),
    .Y(_2298_));
 sky130_fd_sc_hd__nand4_4 _6737_ (.A(_2277_),
    .B(_2284_),
    .C(_2294_),
    .D(_2298_),
    .Y(net88));
 sky130_fd_sc_hd__buf_2 _6738_ (.A(net53),
    .X(_2299_));
 sky130_fd_sc_hd__and2_1 _6739_ (.A(_2007_),
    .B(_2299_),
    .X(_2300_));
 sky130_fd_sc_hd__or2_1 _6740_ (.A(_2007_),
    .B(_2299_),
    .X(_2301_));
 sky130_fd_sc_hd__or2b_1 _6741_ (.A(_2300_),
    .B_N(_2301_),
    .X(_2303_));
 sky130_fd_sc_hd__nor2_1 _6742_ (.A(_1953_),
    .B(_2280_),
    .Y(_2304_));
 sky130_fd_sc_hd__o211ai_1 _6743_ (.A1(_1950_),
    .A2(_1954_),
    .B1(_2279_),
    .C1(_2119_),
    .Y(_2305_));
 sky130_fd_sc_hd__a32o_1 _6744_ (.A1(_1614_),
    .A2(_1955_),
    .A3(_2304_),
    .B1(_2305_),
    .B2(_2278_),
    .X(_2306_));
 sky130_fd_sc_hd__xnor2_1 _6745_ (.A(_2303_),
    .B(_2306_),
    .Y(_2307_));
 sky130_fd_sc_hd__and2b_1 _6746_ (.A_N(_2263_),
    .B(_1821_),
    .X(_2308_));
 sky130_fd_sc_hd__a21o_1 _6747_ (.A1(_2280_),
    .A2(_2296_),
    .B1(_2308_),
    .X(_2309_));
 sky130_fd_sc_hd__or2_1 _6748_ (.A(_2303_),
    .B(_2309_),
    .X(_2310_));
 sky130_fd_sc_hd__nand2_1 _6749_ (.A(_2303_),
    .B(_2309_),
    .Y(_2311_));
 sky130_fd_sc_hd__mux4_1 _6750_ (.A0(_2007_),
    .A1(_1821_),
    .A2(_1810_),
    .A3(_1778_),
    .S0(_0583_),
    .S1(_0584_),
    .X(_2312_));
 sky130_fd_sc_hd__mux2_1 _6751_ (.A0(_1758_),
    .A1(_2312_),
    .S(_0866_),
    .X(_2314_));
 sky130_fd_sc_hd__mux4_1 _6752_ (.A0(_0003_),
    .A1(_0005_),
    .A2(_1018_),
    .A3(_2314_),
    .S0(_0867_),
    .S1(_0573_),
    .X(_2315_));
 sky130_fd_sc_hd__o21ai_1 _6753_ (.A1(_3589_),
    .A2(_2300_),
    .B1(_2301_),
    .Y(_2316_));
 sky130_fd_sc_hd__o22a_1 _6754_ (.A1(_0855_),
    .A2(_2301_),
    .B1(_2316_),
    .B2(_1277_),
    .X(_2317_));
 sky130_fd_sc_hd__a21o_1 _6755_ (.A1(_0854_),
    .A2(_2300_),
    .B1(_2317_),
    .X(_2318_));
 sky130_fd_sc_hd__or2_1 _6756_ (.A(_0783_),
    .B(_3156_),
    .X(_2319_));
 sky130_fd_sc_hd__o31a_1 _6757_ (.A1(_0199_),
    .A2(_0428_),
    .A3(_3163_),
    .B1(_0571_),
    .X(_2320_));
 sky130_fd_sc_hd__a31o_1 _6758_ (.A1(_0573_),
    .A2(_2073_),
    .A3(_3729_),
    .B1(_2320_),
    .X(_2321_));
 sky130_fd_sc_hd__a2bb2o_1 _6759_ (.A1_N(_3730_),
    .A2_N(_2319_),
    .B1(_2321_),
    .B2(_0575_),
    .X(_2322_));
 sky130_fd_sc_hd__a211o_1 _6760_ (.A1(_0844_),
    .A2(_2315_),
    .B1(_2318_),
    .C1(_2322_),
    .X(_2323_));
 sky130_fd_sc_hd__a31o_1 _6761_ (.A1(_3571_),
    .A2(_2310_),
    .A3(_2311_),
    .B1(_2323_),
    .X(_2325_));
 sky130_fd_sc_hd__and2_1 _6762_ (.A(_2128_),
    .B(_2273_),
    .X(_2326_));
 sky130_fd_sc_hd__and2b_1 _6763_ (.A_N(_2271_),
    .B(_2268_),
    .X(_2327_));
 sky130_fd_sc_hd__and2b_1 _6764_ (.A_N(_2131_),
    .B(_2272_),
    .X(_2328_));
 sky130_fd_sc_hd__and2b_1 _6765_ (.A_N(_2265_),
    .B(_2241_),
    .X(_2329_));
 sky130_fd_sc_hd__and2b_1 _6766_ (.A_N(_1982_),
    .B(_2266_),
    .X(_2330_));
 sky130_fd_sc_hd__or2_1 _6767_ (.A(_2238_),
    .B(_2239_),
    .X(_2331_));
 sky130_fd_sc_hd__or2b_1 _6768_ (.A(_2240_),
    .B_N(_2267_),
    .X(_2332_));
 sky130_fd_sc_hd__o211ai_4 _6769_ (.A1(_2011_),
    .A2(_2132_),
    .B1(_2163_),
    .C1(_2164_),
    .Y(_2333_));
 sky130_fd_sc_hd__nor3_1 _6770_ (.A(_2151_),
    .B(_2152_),
    .C(_2162_),
    .Y(_2334_));
 sky130_fd_sc_hd__nand4_2 _6771_ (.A(_0881_),
    .B(_0521_),
    .C(net20),
    .D(net21),
    .Y(_2336_));
 sky130_fd_sc_hd__a22o_1 _6772_ (.A1(_0401_),
    .A2(net20),
    .B1(net21),
    .B2(_0499_),
    .X(_2337_));
 sky130_fd_sc_hd__and2_1 _6773_ (.A(_0303_),
    .B(_1799_),
    .X(_2338_));
 sky130_fd_sc_hd__nand3_1 _6774_ (.A(_2336_),
    .B(_2337_),
    .C(_2338_),
    .Y(_2339_));
 sky130_fd_sc_hd__a21o_1 _6775_ (.A1(_2336_),
    .A2(_2337_),
    .B1(_2338_),
    .X(_2340_));
 sky130_fd_sc_hd__a21bo_1 _6776_ (.A1(_2134_),
    .A2(_2135_),
    .B1_N(_2133_),
    .X(_2341_));
 sky130_fd_sc_hd__nand3_1 _6777_ (.A(_2339_),
    .B(_2340_),
    .C(_2341_),
    .Y(_2342_));
 sky130_fd_sc_hd__a21o_1 _6778_ (.A1(_2339_),
    .A2(_2340_),
    .B1(_2341_),
    .X(_2343_));
 sky130_fd_sc_hd__a22oi_1 _6779_ (.A1(_0052_),
    .A2(_1745_),
    .B1(_1767_),
    .B2(_0183_),
    .Y(_2344_));
 sky130_fd_sc_hd__and4_1 _6780_ (.A(_0172_),
    .B(_0052_),
    .C(_1745_),
    .D(_1767_),
    .X(_2345_));
 sky130_fd_sc_hd__nor2_1 _6781_ (.A(_2344_),
    .B(_2345_),
    .Y(_2347_));
 sky130_fd_sc_hd__nand2_1 _6782_ (.A(_2903_),
    .B(_1952_),
    .Y(_2348_));
 sky130_fd_sc_hd__xnor2_1 _6783_ (.A(_2347_),
    .B(_2348_),
    .Y(_2349_));
 sky130_fd_sc_hd__nand3_1 _6784_ (.A(_2342_),
    .B(_2343_),
    .C(_2349_),
    .Y(_2350_));
 sky130_fd_sc_hd__a21o_1 _6785_ (.A1(_2342_),
    .A2(_2343_),
    .B1(_2349_),
    .X(_2351_));
 sky130_fd_sc_hd__a21bo_1 _6786_ (.A1(_2141_),
    .A2(_2146_),
    .B1_N(_2140_),
    .X(_2352_));
 sky130_fd_sc_hd__and3_2 _6787_ (.A(_2350_),
    .B(_2351_),
    .C(_2352_),
    .X(_2353_));
 sky130_fd_sc_hd__a21oi_1 _6788_ (.A1(_2350_),
    .A2(_2351_),
    .B1(_2352_),
    .Y(_2354_));
 sky130_fd_sc_hd__or2_1 _6789_ (.A(_2155_),
    .B(_2157_),
    .X(_2355_));
 sky130_fd_sc_hd__a32o_1 _6790_ (.A1(_2892_),
    .A2(_1931_),
    .A3(_2143_),
    .B1(_2142_),
    .B2(_1745_),
    .X(_2356_));
 sky130_fd_sc_hd__nand4_2 _6791_ (.A(_3197_),
    .B(_3273_),
    .C(_1898_),
    .D(_1931_),
    .Y(_2358_));
 sky130_fd_sc_hd__a22o_1 _6792_ (.A1(_3272_),
    .A2(_1898_),
    .B1(_1931_),
    .B2(_3197_),
    .X(_2359_));
 sky130_fd_sc_hd__nand4_1 _6793_ (.A(_3386_),
    .B(_1865_),
    .C(_2358_),
    .D(_2359_),
    .Y(_2360_));
 sky130_fd_sc_hd__a22o_1 _6794_ (.A1(_3386_),
    .A2(_1865_),
    .B1(_2358_),
    .B2(_2359_),
    .X(_2361_));
 sky130_fd_sc_hd__and3_1 _6795_ (.A(_2356_),
    .B(_2360_),
    .C(_2361_),
    .X(_2362_));
 sky130_fd_sc_hd__a21o_1 _6796_ (.A1(_2360_),
    .A2(_2361_),
    .B1(_2356_),
    .X(_2363_));
 sky130_fd_sc_hd__and2b_1 _6797_ (.A_N(_2362_),
    .B(_2363_),
    .X(_2364_));
 sky130_fd_sc_hd__xnor2_1 _6798_ (.A(_2355_),
    .B(_2364_),
    .Y(_2365_));
 sky130_fd_sc_hd__or3_1 _6799_ (.A(_2353_),
    .B(_2354_),
    .C(_2365_),
    .X(_2366_));
 sky130_fd_sc_hd__o21ai_1 _6800_ (.A1(_2353_),
    .A2(_2354_),
    .B1(_2365_),
    .Y(_2367_));
 sky130_fd_sc_hd__o211a_1 _6801_ (.A1(_2151_),
    .A2(_2334_),
    .B1(_2366_),
    .C1(_2367_),
    .X(_2369_));
 sky130_fd_sc_hd__a211oi_2 _6802_ (.A1(_2366_),
    .A2(_2367_),
    .B1(_2151_),
    .C1(_2334_),
    .Y(_2370_));
 sky130_fd_sc_hd__or2b_1 _6803_ (.A(_2180_),
    .B_N(_2181_),
    .X(_2371_));
 sky130_fd_sc_hd__or2_1 _6804_ (.A(_2175_),
    .B(_2183_),
    .X(_2372_));
 sky130_fd_sc_hd__or2_1 _6805_ (.A(_2154_),
    .B(_2159_),
    .X(_2373_));
 sky130_fd_sc_hd__nand2_1 _6806_ (.A(_2153_),
    .B(_2161_),
    .Y(_2374_));
 sky130_fd_sc_hd__and4_1 _6807_ (.A(_3720_),
    .B(_0174_),
    .C(_2784_),
    .D(_2510_),
    .X(_2375_));
 sky130_fd_sc_hd__a22o_1 _6808_ (.A1(_0174_),
    .A2(_2784_),
    .B1(_2510_),
    .B2(_3720_),
    .X(_2376_));
 sky130_fd_sc_hd__and4b_1 _6809_ (.A_N(_2375_),
    .B(_0293_),
    .C(_2762_),
    .D(_2376_),
    .X(_2377_));
 sky130_fd_sc_hd__inv_2 _6810_ (.A(_2375_),
    .Y(_2378_));
 sky130_fd_sc_hd__a21boi_1 _6811_ (.A1(_2376_),
    .A2(_2378_),
    .B1_N(_0295_),
    .Y(_2380_));
 sky130_fd_sc_hd__nor2_1 _6812_ (.A(_2377_),
    .B(_2380_),
    .Y(_2381_));
 sky130_fd_sc_hd__and3_1 _6813_ (.A(_3424_),
    .B(_3512_),
    .C(_2576_),
    .X(_2382_));
 sky130_fd_sc_hd__a22o_1 _6814_ (.A1(_3513_),
    .A2(_2576_),
    .B1(_2609_),
    .B2(_3424_),
    .X(_2383_));
 sky130_fd_sc_hd__a21bo_1 _6815_ (.A1(_2609_),
    .A2(_2382_),
    .B1_N(_2383_),
    .X(_2384_));
 sky130_fd_sc_hd__nand2_1 _6816_ (.A(_3685_),
    .B(_2543_),
    .Y(_2385_));
 sky130_fd_sc_hd__xnor2_1 _6817_ (.A(_2384_),
    .B(_2385_),
    .Y(_2386_));
 sky130_fd_sc_hd__a31o_1 _6818_ (.A1(_3685_),
    .A2(_2510_),
    .A3(_2177_),
    .B1(_2176_),
    .X(_2387_));
 sky130_fd_sc_hd__xnor2_1 _6819_ (.A(_2386_),
    .B(_2387_),
    .Y(_2388_));
 sky130_fd_sc_hd__xnor2_1 _6820_ (.A(_2381_),
    .B(_2388_),
    .Y(_2389_));
 sky130_fd_sc_hd__a21oi_1 _6821_ (.A1(_2373_),
    .A2(_2374_),
    .B1(_2389_),
    .Y(_2391_));
 sky130_fd_sc_hd__and3_1 _6822_ (.A(_2373_),
    .B(_2374_),
    .C(_2389_),
    .X(_2392_));
 sky130_fd_sc_hd__a211o_2 _6823_ (.A1(_2371_),
    .A2(_2372_),
    .B1(_2391_),
    .C1(_2392_),
    .X(_2393_));
 sky130_fd_sc_hd__o211ai_2 _6824_ (.A1(_2391_),
    .A2(_2392_),
    .B1(_2371_),
    .C1(_2372_),
    .Y(_2394_));
 sky130_fd_sc_hd__and4bb_2 _6825_ (.A_N(_2369_),
    .B_N(_2370_),
    .C(_2393_),
    .D(_2394_),
    .X(_2395_));
 sky130_fd_sc_hd__a2bb2oi_2 _6826_ (.A1_N(_2369_),
    .A2_N(_2370_),
    .B1(_2393_),
    .B2(_2394_),
    .Y(_2396_));
 sky130_fd_sc_hd__a211oi_4 _6827_ (.A1(_2333_),
    .A2(_2189_),
    .B1(_2395_),
    .C1(_2396_),
    .Y(_2397_));
 sky130_fd_sc_hd__o211a_1 _6828_ (.A1(_2395_),
    .A2(_2396_),
    .B1(_2333_),
    .C1(_2189_),
    .X(_2398_));
 sky130_fd_sc_hd__a21oi_2 _6829_ (.A1(_2214_),
    .A2(_2216_),
    .B1(_2225_),
    .Y(_2399_));
 sky130_fd_sc_hd__a22o_1 _6830_ (.A1(_2456_),
    .A2(_1170_),
    .B1(_1295_),
    .B2(_2390_),
    .X(_2400_));
 sky130_fd_sc_hd__and4_1 _6831_ (.A(_2390_),
    .B(_2456_),
    .C(_1169_),
    .D(_1294_),
    .X(_2402_));
 sky130_fd_sc_hd__inv_2 _6832_ (.A(_2402_),
    .Y(_2403_));
 sky130_fd_sc_hd__a22oi_1 _6833_ (.A1(_2335_),
    .A2(_1448_),
    .B1(_2400_),
    .B2(_2403_),
    .Y(_2404_));
 sky130_fd_sc_hd__and4b_1 _6834_ (.A_N(_2402_),
    .B(_1448_),
    .C(_2335_),
    .D(_2400_),
    .X(_2405_));
 sky130_fd_sc_hd__or2_1 _6835_ (.A(_2404_),
    .B(_2405_),
    .X(_2406_));
 sky130_fd_sc_hd__a22o_1 _6836_ (.A1(_2226_),
    .A2(_0721_),
    .B1(_0874_),
    .B2(_2171_),
    .X(_2407_));
 sky130_fd_sc_hd__nand4_1 _6837_ (.A(_2171_),
    .B(_2226_),
    .C(_0721_),
    .D(_0874_),
    .Y(_2408_));
 sky130_fd_sc_hd__a22oi_1 _6838_ (.A1(_2127_),
    .A2(_1008_),
    .B1(_2407_),
    .B2(_2408_),
    .Y(_2409_));
 sky130_fd_sc_hd__and4_1 _6839_ (.A(_2127_),
    .B(_1007_),
    .C(_2407_),
    .D(_2408_),
    .X(_2410_));
 sky130_fd_sc_hd__a21bo_1 _6840_ (.A1(_2205_),
    .A2(_2207_),
    .B1_N(_2203_),
    .X(_2411_));
 sky130_fd_sc_hd__or3b_2 _6841_ (.A(_2409_),
    .B(_2410_),
    .C_N(_2411_),
    .X(_2413_));
 sky130_fd_sc_hd__o21bai_1 _6842_ (.A1(_2409_),
    .A2(_2410_),
    .B1_N(_2411_),
    .Y(_2414_));
 sky130_fd_sc_hd__nand2_1 _6843_ (.A(_2413_),
    .B(_2414_),
    .Y(_2415_));
 sky130_fd_sc_hd__or2_2 _6844_ (.A(_2406_),
    .B(_2415_),
    .X(_2416_));
 sky130_fd_sc_hd__nand2_1 _6845_ (.A(_2406_),
    .B(_2415_),
    .Y(_2417_));
 sky130_fd_sc_hd__and2_1 _6846_ (.A(_2416_),
    .B(_2417_),
    .X(_2418_));
 sky130_fd_sc_hd__or2_1 _6847_ (.A(_2218_),
    .B(_2223_),
    .X(_2419_));
 sky130_fd_sc_hd__nand2_1 _6848_ (.A(_2217_),
    .B(_2224_),
    .Y(_2420_));
 sky130_fd_sc_hd__or2_1 _6849_ (.A(_2219_),
    .B(_2221_),
    .X(_2421_));
 sky130_fd_sc_hd__a22o_1 _6850_ (.A1(_2707_),
    .A2(_0327_),
    .B1(_0454_),
    .B2(_2664_),
    .X(_2422_));
 sky130_fd_sc_hd__nand4_1 _6851_ (.A(_2664_),
    .B(_2718_),
    .C(_0328_),
    .D(_0454_),
    .Y(_2424_));
 sky130_fd_sc_hd__a22oi_2 _6852_ (.A1(_2270_),
    .A2(_0689_),
    .B1(_2422_),
    .B2(_2424_),
    .Y(_2425_));
 sky130_fd_sc_hd__and4_1 _6853_ (.A(_2270_),
    .B(_0688_),
    .C(_2422_),
    .D(_2424_),
    .X(_2426_));
 sky130_fd_sc_hd__a211o_1 _6854_ (.A1(_2172_),
    .A2(_2174_),
    .B1(_2425_),
    .C1(_2426_),
    .X(_2427_));
 sky130_fd_sc_hd__o211ai_1 _6855_ (.A1(_2425_),
    .A2(_2426_),
    .B1(_2172_),
    .C1(_2174_),
    .Y(_2428_));
 sky130_fd_sc_hd__and2_1 _6856_ (.A(_2427_),
    .B(_2428_),
    .X(_2429_));
 sky130_fd_sc_hd__xnor2_1 _6857_ (.A(_2421_),
    .B(_2429_),
    .Y(_2430_));
 sky130_fd_sc_hd__a21o_1 _6858_ (.A1(_2419_),
    .A2(_2420_),
    .B1(_2430_),
    .X(_2431_));
 sky130_fd_sc_hd__nand3_1 _6859_ (.A(_2419_),
    .B(_2420_),
    .C(_2430_),
    .Y(_2432_));
 sky130_fd_sc_hd__nand3_2 _6860_ (.A(_2418_),
    .B(_2431_),
    .C(_2432_),
    .Y(_2433_));
 sky130_fd_sc_hd__a21o_1 _6861_ (.A1(_2431_),
    .A2(_2432_),
    .B1(_2418_),
    .X(_2435_));
 sky130_fd_sc_hd__o211ai_4 _6862_ (.A1(_2185_),
    .A2(_2187_),
    .B1(_2433_),
    .C1(_2435_),
    .Y(_2436_));
 sky130_fd_sc_hd__a211o_1 _6863_ (.A1(_2433_),
    .A2(_2435_),
    .B1(_2185_),
    .C1(_2187_),
    .X(_2437_));
 sky130_fd_sc_hd__o211ai_4 _6864_ (.A1(_2399_),
    .A2(_2229_),
    .B1(_2436_),
    .C1(_2437_),
    .Y(_2438_));
 sky130_fd_sc_hd__a211o_1 _6865_ (.A1(_2436_),
    .A2(_2437_),
    .B1(_2399_),
    .C1(_2229_),
    .X(_2439_));
 sky130_fd_sc_hd__and4bb_2 _6866_ (.A_N(_2397_),
    .B_N(_2398_),
    .C(_2438_),
    .D(_2439_),
    .X(_2440_));
 sky130_fd_sc_hd__a2bb2o_1 _6867_ (.A1_N(_2397_),
    .A2_N(_2398_),
    .B1(_2438_),
    .B2(_2439_),
    .X(_2441_));
 sky130_fd_sc_hd__and2b_1 _6868_ (.A_N(_2440_),
    .B(_2441_),
    .X(_2442_));
 sky130_fd_sc_hd__nor2_1 _6869_ (.A(_2191_),
    .B(_2235_),
    .Y(_2443_));
 sky130_fd_sc_hd__xnor2_1 _6870_ (.A(_2442_),
    .B(_2443_),
    .Y(_2444_));
 sky130_fd_sc_hd__or2_1 _6871_ (.A(_2258_),
    .B(_2261_),
    .X(_2446_));
 sky130_fd_sc_hd__nand3_1 _6872_ (.A(_3209_),
    .B(_2263_),
    .C(_2262_),
    .Y(_2447_));
 sky130_fd_sc_hd__a22oi_2 _6873_ (.A1(_1067_),
    .A2(_2263_),
    .B1(_2299_),
    .B2(_3209_),
    .Y(_2448_));
 sky130_fd_sc_hd__and4_2 _6874_ (.A(_1067_),
    .B(_1384_),
    .C(_2263_),
    .D(_2299_),
    .X(_2449_));
 sky130_fd_sc_hd__and2b_1 _6875_ (.A_N(_2254_),
    .B(_2243_),
    .X(_2450_));
 sky130_fd_sc_hd__inv_2 _6876_ (.A(_2450_),
    .Y(_2451_));
 sky130_fd_sc_hd__or2_1 _6877_ (.A(_2255_),
    .B(_2257_),
    .X(_2452_));
 sky130_fd_sc_hd__or2b_1 _6878_ (.A(_2252_),
    .B_N(_2245_),
    .X(_2453_));
 sky130_fd_sc_hd__nand2_1 _6879_ (.A(_2244_),
    .B(_2253_),
    .Y(_2454_));
 sky130_fd_sc_hd__or2b_1 _6880_ (.A(_2208_),
    .B_N(_2209_),
    .X(_2455_));
 sky130_fd_sc_hd__or2_1 _6881_ (.A(_2249_),
    .B(_2251_),
    .X(_2457_));
 sky130_fd_sc_hd__a22oi_1 _6882_ (.A1(_0106_),
    .A2(_1607_),
    .B1(net50),
    .B2(_0215_),
    .Y(_2458_));
 sky130_fd_sc_hd__and4_1 _6883_ (.A(_0106_),
    .B(_0215_),
    .C(_1607_),
    .D(net50),
    .X(_2459_));
 sky130_fd_sc_hd__o2bb2a_1 _6884_ (.A1_N(_0357_),
    .A2_N(_1949_),
    .B1(_2458_),
    .B2(_2459_),
    .X(_2460_));
 sky130_fd_sc_hd__and4bb_1 _6885_ (.A_N(_2458_),
    .B_N(_2459_),
    .C(_0357_),
    .D(_1949_),
    .X(_2461_));
 sky130_fd_sc_hd__a211o_1 _6886_ (.A1(_2199_),
    .A2(_2201_),
    .B1(_2460_),
    .C1(_2461_),
    .X(_2462_));
 sky130_fd_sc_hd__o211ai_1 _6887_ (.A1(_2460_),
    .A2(_2461_),
    .B1(_2199_),
    .C1(_2201_),
    .Y(_2463_));
 sky130_fd_sc_hd__and2_1 _6888_ (.A(_2462_),
    .B(_2463_),
    .X(_2464_));
 sky130_fd_sc_hd__xnor2_1 _6889_ (.A(_2457_),
    .B(_2464_),
    .Y(_2465_));
 sky130_fd_sc_hd__a21oi_2 _6890_ (.A1(_2455_),
    .A2(_2211_),
    .B1(_2465_),
    .Y(_2466_));
 sky130_fd_sc_hd__and3_1 _6891_ (.A(_2455_),
    .B(_2211_),
    .C(_2465_),
    .X(_2468_));
 sky130_fd_sc_hd__a211oi_2 _6892_ (.A1(_2453_),
    .A2(_2454_),
    .B1(_2466_),
    .C1(_2468_),
    .Y(_2469_));
 sky130_fd_sc_hd__o211a_1 _6893_ (.A1(_2466_),
    .A2(_2468_),
    .B1(_2453_),
    .C1(_2454_),
    .X(_2470_));
 sky130_fd_sc_hd__a211oi_2 _6894_ (.A1(_2451_),
    .A2(_2452_),
    .B1(_2469_),
    .C1(_2470_),
    .Y(_2471_));
 sky130_fd_sc_hd__o211a_1 _6895_ (.A1(_2469_),
    .A2(_2470_),
    .B1(_2451_),
    .C1(_2452_),
    .X(_2472_));
 sky130_fd_sc_hd__nor4_1 _6896_ (.A(_2448_),
    .B(_2449_),
    .C(_2471_),
    .D(_2472_),
    .Y(_2473_));
 sky130_fd_sc_hd__o22a_1 _6897_ (.A1(_2448_),
    .A2(_2449_),
    .B1(_2471_),
    .B2(_2472_),
    .X(_2474_));
 sky130_fd_sc_hd__a211o_1 _6898_ (.A1(_2231_),
    .A2(_2233_),
    .B1(_2473_),
    .C1(_2474_),
    .X(_2475_));
 sky130_fd_sc_hd__inv_2 _6899_ (.A(_2475_),
    .Y(_2476_));
 sky130_fd_sc_hd__o211a_1 _6900_ (.A1(_2473_),
    .A2(_2474_),
    .B1(_2231_),
    .C1(_2233_),
    .X(_2477_));
 sky130_fd_sc_hd__a211o_1 _6901_ (.A1(_2446_),
    .A2(_2447_),
    .B1(_2476_),
    .C1(_2477_),
    .X(_2479_));
 sky130_fd_sc_hd__o211ai_1 _6902_ (.A1(_2476_),
    .A2(_2477_),
    .B1(_2446_),
    .C1(_2447_),
    .Y(_2480_));
 sky130_fd_sc_hd__and3_2 _6903_ (.A(_2444_),
    .B(_2479_),
    .C(_2480_),
    .X(_2481_));
 sky130_fd_sc_hd__a21oi_1 _6904_ (.A1(_2479_),
    .A2(_2480_),
    .B1(_2444_),
    .Y(_2482_));
 sky130_fd_sc_hd__a211o_2 _6905_ (.A1(_2331_),
    .A2(_2332_),
    .B1(_2481_),
    .C1(_2482_),
    .X(_2483_));
 sky130_fd_sc_hd__o211ai_2 _6906_ (.A1(_2481_),
    .A2(_2482_),
    .B1(_2331_),
    .C1(_2332_),
    .Y(_2484_));
 sky130_fd_sc_hd__o211ai_4 _6907_ (.A1(_2329_),
    .A2(_2330_),
    .B1(_2483_),
    .C1(_2484_),
    .Y(_2485_));
 sky130_fd_sc_hd__a211o_1 _6908_ (.A1(_2483_),
    .A2(_2484_),
    .B1(_2329_),
    .C1(_2330_),
    .X(_2486_));
 sky130_fd_sc_hd__o211ai_4 _6909_ (.A1(_2327_),
    .A2(_2328_),
    .B1(_2485_),
    .C1(_2486_),
    .Y(_2487_));
 sky130_fd_sc_hd__a211o_1 _6910_ (.A1(_2485_),
    .A2(_2486_),
    .B1(_2327_),
    .C1(_2328_),
    .X(_2488_));
 sky130_fd_sc_hd__and2_1 _6911_ (.A(_2487_),
    .B(_2488_),
    .X(_2490_));
 sky130_fd_sc_hd__xor2_1 _6912_ (.A(_2326_),
    .B(_2490_),
    .X(_2491_));
 sky130_fd_sc_hd__or4_1 _6913_ (.A(_1754_),
    .B(_1926_),
    .C(_2105_),
    .D(_2275_),
    .X(_2492_));
 sky130_fd_sc_hd__a31oi_1 _6914_ (.A1(net129),
    .A2(_1620_),
    .A3(_1623_),
    .B1(_2492_),
    .Y(_2493_));
 sky130_fd_sc_hd__nor3_1 _6915_ (.A(_2105_),
    .B(_2107_),
    .C(_2275_),
    .Y(_2494_));
 sky130_fd_sc_hd__a21oi_1 _6916_ (.A1(_2102_),
    .A2(_2126_),
    .B1(_2274_),
    .Y(_2495_));
 sky130_fd_sc_hd__or4_1 _6917_ (.A(_2491_),
    .B(_2493_),
    .C(_2494_),
    .D(_2495_),
    .X(_2496_));
 sky130_fd_sc_hd__o31ai_2 _6918_ (.A1(net168),
    .A2(_2494_),
    .A3(_2495_),
    .B1(_2491_),
    .Y(_2497_));
 sky130_fd_sc_hd__and3_1 _6919_ (.A(_0320_),
    .B(_2496_),
    .C(_2497_),
    .X(_2498_));
 sky130_fd_sc_hd__a211o_1 _6920_ (.A1(_0419_),
    .A2(_2307_),
    .B1(_2325_),
    .C1(_2498_),
    .X(net89));
 sky130_fd_sc_hd__nand2_1 _6921_ (.A(_2326_),
    .B(_2490_),
    .Y(_2500_));
 sky130_fd_sc_hd__inv_2 _6922_ (.A(_2487_),
    .Y(_2501_));
 sky130_fd_sc_hd__and2b_1 _6923_ (.A_N(_2443_),
    .B(_2442_),
    .X(_2502_));
 sky130_fd_sc_hd__nor3_1 _6924_ (.A(_2353_),
    .B(_2354_),
    .C(_2365_),
    .Y(_2503_));
 sky130_fd_sc_hd__a22o_1 _6925_ (.A1(_0521_),
    .A2(net21),
    .B1(net22),
    .B2(_0881_),
    .X(_2504_));
 sky130_fd_sc_hd__nand4_2 _6926_ (.A(_0881_),
    .B(_0521_),
    .C(net21),
    .D(net22),
    .Y(_2505_));
 sky130_fd_sc_hd__and2_1 _6927_ (.A(_0303_),
    .B(net20),
    .X(_2506_));
 sky130_fd_sc_hd__a21o_1 _6928_ (.A1(_2504_),
    .A2(_2505_),
    .B1(_2506_),
    .X(_2507_));
 sky130_fd_sc_hd__nand3_1 _6929_ (.A(_2504_),
    .B(_2505_),
    .C(_2506_),
    .Y(_2508_));
 sky130_fd_sc_hd__a21bo_1 _6930_ (.A1(_2337_),
    .A2(_2338_),
    .B1_N(_2336_),
    .X(_2509_));
 sky130_fd_sc_hd__nand3_1 _6931_ (.A(_2507_),
    .B(_2508_),
    .C(_2509_),
    .Y(_2511_));
 sky130_fd_sc_hd__a21o_1 _6932_ (.A1(_2507_),
    .A2(_2508_),
    .B1(_2509_),
    .X(_2512_));
 sky130_fd_sc_hd__a22oi_1 _6933_ (.A1(_0052_),
    .A2(_1767_),
    .B1(_1799_),
    .B2(_0183_),
    .Y(_2513_));
 sky130_fd_sc_hd__and4_1 _6934_ (.A(_0172_),
    .B(_0052_),
    .C(_1767_),
    .D(_1799_),
    .X(_2514_));
 sky130_fd_sc_hd__nor2_1 _6935_ (.A(_2513_),
    .B(_2514_),
    .Y(_2515_));
 sky130_fd_sc_hd__nand2_1 _6936_ (.A(_2903_),
    .B(_1745_),
    .Y(_2516_));
 sky130_fd_sc_hd__xnor2_1 _6937_ (.A(_2515_),
    .B(_2516_),
    .Y(_2517_));
 sky130_fd_sc_hd__nand3_1 _6938_ (.A(_2511_),
    .B(_2512_),
    .C(_2517_),
    .Y(_2518_));
 sky130_fd_sc_hd__a21o_1 _6939_ (.A1(_2511_),
    .A2(_2512_),
    .B1(_2517_),
    .X(_2519_));
 sky130_fd_sc_hd__a21bo_1 _6940_ (.A1(_2343_),
    .A2(_2349_),
    .B1_N(_2342_),
    .X(_2520_));
 sky130_fd_sc_hd__and3_2 _6941_ (.A(_2518_),
    .B(_2519_),
    .C(_2520_),
    .X(_2522_));
 sky130_fd_sc_hd__a21oi_2 _6942_ (.A1(_2518_),
    .A2(_2519_),
    .B1(_2520_),
    .Y(_2523_));
 sky130_fd_sc_hd__nand2_1 _6943_ (.A(_2358_),
    .B(_2360_),
    .Y(_2524_));
 sky130_fd_sc_hd__a31o_1 _6944_ (.A1(_2903_),
    .A2(_1952_),
    .A3(_2347_),
    .B1(_2345_),
    .X(_2525_));
 sky130_fd_sc_hd__a22oi_1 _6945_ (.A1(_3273_),
    .A2(_1931_),
    .B1(_1952_),
    .B2(_3198_),
    .Y(_2526_));
 sky130_fd_sc_hd__and4_1 _6946_ (.A(_3197_),
    .B(_3273_),
    .C(_1931_),
    .D(_1952_),
    .X(_2527_));
 sky130_fd_sc_hd__nor2_1 _6947_ (.A(_2526_),
    .B(_2527_),
    .Y(_2528_));
 sky130_fd_sc_hd__nand2_1 _6948_ (.A(_3386_),
    .B(_1898_),
    .Y(_2529_));
 sky130_fd_sc_hd__xnor2_2 _6949_ (.A(_2528_),
    .B(_2529_),
    .Y(_2530_));
 sky130_fd_sc_hd__xor2_2 _6950_ (.A(_2525_),
    .B(_2530_),
    .X(_2531_));
 sky130_fd_sc_hd__xnor2_2 _6951_ (.A(_2524_),
    .B(_2531_),
    .Y(_2533_));
 sky130_fd_sc_hd__or3_1 _6952_ (.A(_2522_),
    .B(_2523_),
    .C(_2533_),
    .X(_2534_));
 sky130_fd_sc_hd__o21ai_2 _6953_ (.A1(_2522_),
    .A2(_2523_),
    .B1(_2533_),
    .Y(_2535_));
 sky130_fd_sc_hd__o211ai_2 _6954_ (.A1(_2353_),
    .A2(_2503_),
    .B1(_2534_),
    .C1(_2535_),
    .Y(_2536_));
 sky130_fd_sc_hd__a211o_1 _6955_ (.A1(_2534_),
    .A2(_2535_),
    .B1(_2353_),
    .C1(_2503_),
    .X(_2537_));
 sky130_fd_sc_hd__or2b_1 _6956_ (.A(_2387_),
    .B_N(_2386_),
    .X(_2538_));
 sky130_fd_sc_hd__and2b_1 _6957_ (.A_N(_2386_),
    .B(_2387_),
    .X(_2539_));
 sky130_fd_sc_hd__a21oi_1 _6958_ (.A1(_2381_),
    .A2(_2538_),
    .B1(_2539_),
    .Y(_2540_));
 sky130_fd_sc_hd__a21o_1 _6959_ (.A1(_2355_),
    .A2(_2363_),
    .B1(_2362_),
    .X(_2541_));
 sky130_fd_sc_hd__and3_1 _6960_ (.A(_3719_),
    .B(_0100_),
    .C(_2499_),
    .X(_2542_));
 sky130_fd_sc_hd__a22o_1 _6961_ (.A1(_0100_),
    .A2(_2499_),
    .B1(_2543_),
    .B2(_3719_),
    .X(_2544_));
 sky130_fd_sc_hd__a21bo_1 _6962_ (.A1(_2543_),
    .A2(_2542_),
    .B1_N(_2544_),
    .X(_2545_));
 sky130_fd_sc_hd__nand2_1 _6963_ (.A(_0293_),
    .B(_2784_),
    .Y(_2546_));
 sky130_fd_sc_hd__xor2_2 _6964_ (.A(_2545_),
    .B(_2546_),
    .X(_2547_));
 sky130_fd_sc_hd__a22o_1 _6965_ (.A1(_3513_),
    .A2(_2609_),
    .B1(_1865_),
    .B2(_3424_),
    .X(_2548_));
 sky130_fd_sc_hd__nand4_4 _6966_ (.A(_3424_),
    .B(_3513_),
    .C(_2609_),
    .D(_1865_),
    .Y(_2549_));
 sky130_fd_sc_hd__a22o_1 _6967_ (.A1(_3685_),
    .A2(_2576_),
    .B1(_2548_),
    .B2(_2549_),
    .X(_2550_));
 sky130_fd_sc_hd__nand4_4 _6968_ (.A(_3685_),
    .B(_2576_),
    .C(_2548_),
    .D(_2549_),
    .Y(_2551_));
 sky130_fd_sc_hd__a32o_1 _6969_ (.A1(_3620_),
    .A2(_2543_),
    .A3(_2383_),
    .B1(_2382_),
    .B2(_2609_),
    .X(_2552_));
 sky130_fd_sc_hd__nand3_4 _6970_ (.A(_2550_),
    .B(_2551_),
    .C(_2552_),
    .Y(_2553_));
 sky130_fd_sc_hd__a21o_1 _6971_ (.A1(_2550_),
    .A2(_2551_),
    .B1(_2552_),
    .X(_2555_));
 sky130_fd_sc_hd__nand3_4 _6972_ (.A(_2547_),
    .B(_2553_),
    .C(_2555_),
    .Y(_2556_));
 sky130_fd_sc_hd__a21o_1 _6973_ (.A1(_2553_),
    .A2(_2555_),
    .B1(_2547_),
    .X(_2557_));
 sky130_fd_sc_hd__and3_1 _6974_ (.A(_2541_),
    .B(_2556_),
    .C(_2557_),
    .X(_2558_));
 sky130_fd_sc_hd__a21oi_1 _6975_ (.A1(_2556_),
    .A2(_2557_),
    .B1(_2541_),
    .Y(_2559_));
 sky130_fd_sc_hd__or3_2 _6976_ (.A(_2540_),
    .B(_2558_),
    .C(_2559_),
    .X(_2560_));
 sky130_fd_sc_hd__o21ai_2 _6977_ (.A1(_2558_),
    .A2(_2559_),
    .B1(_2540_),
    .Y(_2561_));
 sky130_fd_sc_hd__nand4_2 _6978_ (.A(_2536_),
    .B(_2537_),
    .C(_2560_),
    .D(_2561_),
    .Y(_2562_));
 sky130_fd_sc_hd__a22o_1 _6979_ (.A1(_2536_),
    .A2(_2537_),
    .B1(_2560_),
    .B2(_2561_),
    .X(_2563_));
 sky130_fd_sc_hd__o211a_1 _6980_ (.A1(_2369_),
    .A2(_2395_),
    .B1(_2562_),
    .C1(_2563_),
    .X(_2564_));
 sky130_fd_sc_hd__a211oi_2 _6981_ (.A1(_2562_),
    .A2(_2563_),
    .B1(_2369_),
    .C1(_2395_),
    .Y(_2566_));
 sky130_fd_sc_hd__inv_2 _6982_ (.A(_2431_),
    .Y(_2567_));
 sky130_fd_sc_hd__and3_1 _6983_ (.A(_2418_),
    .B(_2431_),
    .C(_2432_),
    .X(_2568_));
 sky130_fd_sc_hd__a21o_1 _6984_ (.A1(_2373_),
    .A2(_2374_),
    .B1(_2389_),
    .X(_2569_));
 sky130_fd_sc_hd__a22o_1 _6985_ (.A1(_2127_),
    .A2(_1169_),
    .B1(_1294_),
    .B2(_2456_),
    .X(_2570_));
 sky130_fd_sc_hd__inv_2 _6986_ (.A(_2570_),
    .Y(_2571_));
 sky130_fd_sc_hd__and4_1 _6987_ (.A(_2456_),
    .B(_2127_),
    .C(_1169_),
    .D(_1295_),
    .X(_2572_));
 sky130_fd_sc_hd__o2bb2a_1 _6988_ (.A1_N(_2401_),
    .A2_N(_1448_),
    .B1(_2571_),
    .B2(_2572_),
    .X(_2573_));
 sky130_fd_sc_hd__and4b_1 _6989_ (.A_N(_2572_),
    .B(net48),
    .C(_2401_),
    .D(_2570_),
    .X(_2574_));
 sky130_fd_sc_hd__or2_1 _6990_ (.A(_2573_),
    .B(_2574_),
    .X(_2575_));
 sky130_fd_sc_hd__a22oi_1 _6991_ (.A1(_2270_),
    .A2(_0722_),
    .B1(_0875_),
    .B2(_2226_),
    .Y(_2577_));
 sky130_fd_sc_hd__and4_1 _6992_ (.A(_2226_),
    .B(_2270_),
    .C(_0721_),
    .D(_0874_),
    .X(_2578_));
 sky130_fd_sc_hd__o2bb2a_1 _6993_ (.A1_N(_2171_),
    .A2_N(_1008_),
    .B1(_2577_),
    .B2(_2578_),
    .X(_2579_));
 sky130_fd_sc_hd__and4bb_1 _6994_ (.A_N(_2577_),
    .B_N(_2578_),
    .C(_2171_),
    .D(_1008_),
    .X(_2580_));
 sky130_fd_sc_hd__nor2_1 _6995_ (.A(_2579_),
    .B(_2580_),
    .Y(_2581_));
 sky130_fd_sc_hd__a41o_1 _6996_ (.A1(_2171_),
    .A2(_2226_),
    .A3(_0722_),
    .A4(_0875_),
    .B1(_2410_),
    .X(_2582_));
 sky130_fd_sc_hd__xnor2_1 _6997_ (.A(_2581_),
    .B(_2582_),
    .Y(_2583_));
 sky130_fd_sc_hd__or2_1 _6998_ (.A(_2575_),
    .B(_2583_),
    .X(_2584_));
 sky130_fd_sc_hd__nand2_1 _6999_ (.A(_2575_),
    .B(_2583_),
    .Y(_2585_));
 sky130_fd_sc_hd__and2_1 _7000_ (.A(_2584_),
    .B(_2585_),
    .X(_2586_));
 sky130_fd_sc_hd__nand2_1 _7001_ (.A(_2421_),
    .B(_2429_),
    .Y(_2588_));
 sky130_fd_sc_hd__a41o_1 _7002_ (.A1(_2675_),
    .A2(_2718_),
    .A3(_0328_),
    .A4(_0559_),
    .B1(_2426_),
    .X(_2589_));
 sky130_fd_sc_hd__a22o_1 _7003_ (.A1(_2762_),
    .A2(_0328_),
    .B1(_0559_),
    .B2(_2718_),
    .X(_2590_));
 sky130_fd_sc_hd__nand4_2 _7004_ (.A(_2718_),
    .B(_2762_),
    .C(_0328_),
    .D(_0559_),
    .Y(_2591_));
 sky130_fd_sc_hd__a22o_1 _7005_ (.A1(_2664_),
    .A2(_0689_),
    .B1(_2590_),
    .B2(_2591_),
    .X(_2592_));
 sky130_fd_sc_hd__nand4_2 _7006_ (.A(_2664_),
    .B(_0689_),
    .C(_2590_),
    .D(_2591_),
    .Y(_2593_));
 sky130_fd_sc_hd__o211ai_1 _7007_ (.A1(_2375_),
    .A2(_2377_),
    .B1(_2592_),
    .C1(_2593_),
    .Y(_2594_));
 sky130_fd_sc_hd__a211o_1 _7008_ (.A1(_2592_),
    .A2(_2593_),
    .B1(_2375_),
    .C1(_2377_),
    .X(_2595_));
 sky130_fd_sc_hd__nand2_1 _7009_ (.A(_2594_),
    .B(_2595_),
    .Y(_2596_));
 sky130_fd_sc_hd__xor2_1 _7010_ (.A(_2589_),
    .B(_2596_),
    .X(_2597_));
 sky130_fd_sc_hd__a21o_1 _7011_ (.A1(_2427_),
    .A2(_2588_),
    .B1(_2597_),
    .X(_2599_));
 sky130_fd_sc_hd__nand3_2 _7012_ (.A(_2427_),
    .B(_2588_),
    .C(_2597_),
    .Y(_2600_));
 sky130_fd_sc_hd__and3_1 _7013_ (.A(_2586_),
    .B(_2599_),
    .C(_2600_),
    .X(_2601_));
 sky130_fd_sc_hd__a21oi_2 _7014_ (.A1(_2599_),
    .A2(_2600_),
    .B1(_2586_),
    .Y(_2602_));
 sky130_fd_sc_hd__a211o_2 _7015_ (.A1(_2569_),
    .A2(_2393_),
    .B1(_2601_),
    .C1(_2602_),
    .X(_2603_));
 sky130_fd_sc_hd__o211ai_4 _7016_ (.A1(_2601_),
    .A2(_2602_),
    .B1(_2569_),
    .C1(_2393_),
    .Y(_2604_));
 sky130_fd_sc_hd__o211ai_4 _7017_ (.A1(_2567_),
    .A2(_2568_),
    .B1(_2603_),
    .C1(_2604_),
    .Y(_2605_));
 sky130_fd_sc_hd__a211o_1 _7018_ (.A1(_2603_),
    .A2(_2604_),
    .B1(_2567_),
    .C1(_2568_),
    .X(_2606_));
 sky130_fd_sc_hd__or4bb_2 _7019_ (.A(_2564_),
    .B(_2566_),
    .C_N(_2605_),
    .D_N(_2606_),
    .X(_2607_));
 sky130_fd_sc_hd__a2bb2o_1 _7020_ (.A1_N(_2564_),
    .A2_N(_2566_),
    .B1(_2605_),
    .B2(_2606_),
    .X(_2608_));
 sky130_fd_sc_hd__o211ai_4 _7021_ (.A1(_2397_),
    .A2(_2440_),
    .B1(_2607_),
    .C1(_2608_),
    .Y(_2610_));
 sky130_fd_sc_hd__a211o_1 _7022_ (.A1(_2607_),
    .A2(_2608_),
    .B1(_2397_),
    .C1(_2440_),
    .X(_2611_));
 sky130_fd_sc_hd__inv_2 _7023_ (.A(_2471_),
    .Y(_2612_));
 sky130_fd_sc_hd__or4_1 _7024_ (.A(_2448_),
    .B(_2449_),
    .C(_2471_),
    .D(_2472_),
    .X(_2613_));
 sky130_fd_sc_hd__inv_2 _7025_ (.A(_2449_),
    .Y(_2614_));
 sky130_fd_sc_hd__a22o_1 _7026_ (.A1(_1045_),
    .A2(net52),
    .B1(_2299_),
    .B2(_1056_),
    .X(_2615_));
 sky130_fd_sc_hd__inv_2 _7027_ (.A(_2615_),
    .Y(_2616_));
 sky130_fd_sc_hd__and4_1 _7028_ (.A(_0357_),
    .B(_1056_),
    .C(net52),
    .D(net53),
    .X(_2617_));
 sky130_fd_sc_hd__o2bb2a_1 _7029_ (.A1_N(_1384_),
    .A2_N(net54),
    .B1(_2616_),
    .B2(_2617_),
    .X(_2618_));
 sky130_fd_sc_hd__and4b_1 _7030_ (.A_N(_2617_),
    .B(net54),
    .C(_1002_),
    .D(_2615_),
    .X(_2619_));
 sky130_fd_sc_hd__or2_1 _7031_ (.A(_2618_),
    .B(_2619_),
    .X(_2621_));
 sky130_fd_sc_hd__nor2_1 _7032_ (.A(_2614_),
    .B(_2621_),
    .Y(_2622_));
 sky130_fd_sc_hd__and2_1 _7033_ (.A(_2614_),
    .B(_2621_),
    .X(_2623_));
 sky130_fd_sc_hd__or2_1 _7034_ (.A(_2622_),
    .B(_2623_),
    .X(_2624_));
 sky130_fd_sc_hd__inv_2 _7035_ (.A(_2466_),
    .Y(_2625_));
 sky130_fd_sc_hd__a211o_1 _7036_ (.A1(_2453_),
    .A2(_2454_),
    .B1(_2466_),
    .C1(_2468_),
    .X(_2626_));
 sky130_fd_sc_hd__nand2_1 _7037_ (.A(_2457_),
    .B(_2464_),
    .Y(_2627_));
 sky130_fd_sc_hd__or2_2 _7038_ (.A(_2459_),
    .B(_2461_),
    .X(_2628_));
 sky130_fd_sc_hd__or2_1 _7039_ (.A(_2402_),
    .B(_2405_),
    .X(_2629_));
 sky130_fd_sc_hd__a22o_1 _7040_ (.A1(_2335_),
    .A2(_1607_),
    .B1(_1797_),
    .B2(_0117_),
    .X(_2630_));
 sky130_fd_sc_hd__nand4_1 _7041_ (.A(_0117_),
    .B(_2335_),
    .C(_1607_),
    .D(_1797_),
    .Y(_2632_));
 sky130_fd_sc_hd__a22oi_1 _7042_ (.A1(_0226_),
    .A2(_1949_),
    .B1(_2630_),
    .B2(_2632_),
    .Y(_2633_));
 sky130_fd_sc_hd__and4_1 _7043_ (.A(_0226_),
    .B(_1949_),
    .C(_2630_),
    .D(_2632_),
    .X(_2634_));
 sky130_fd_sc_hd__or2_1 _7044_ (.A(_2633_),
    .B(_2634_),
    .X(_2635_));
 sky130_fd_sc_hd__xnor2_2 _7045_ (.A(_2629_),
    .B(_2635_),
    .Y(_2636_));
 sky130_fd_sc_hd__xnor2_2 _7046_ (.A(_2628_),
    .B(_2636_),
    .Y(_2637_));
 sky130_fd_sc_hd__a21oi_4 _7047_ (.A1(_2413_),
    .A2(_2416_),
    .B1(_2637_),
    .Y(_2638_));
 sky130_fd_sc_hd__and3_1 _7048_ (.A(_2413_),
    .B(_2416_),
    .C(_2637_),
    .X(_2639_));
 sky130_fd_sc_hd__a211oi_4 _7049_ (.A1(_2462_),
    .A2(_2627_),
    .B1(_2638_),
    .C1(_2639_),
    .Y(_2640_));
 sky130_fd_sc_hd__o211a_1 _7050_ (.A1(_2638_),
    .A2(_2639_),
    .B1(_2462_),
    .C1(_2627_),
    .X(_2641_));
 sky130_fd_sc_hd__a211oi_2 _7051_ (.A1(_2625_),
    .A2(_2626_),
    .B1(_2640_),
    .C1(_2641_),
    .Y(_2643_));
 sky130_fd_sc_hd__o211a_1 _7052_ (.A1(_2640_),
    .A2(_2641_),
    .B1(_2625_),
    .C1(_2626_),
    .X(_2644_));
 sky130_fd_sc_hd__nor3_1 _7053_ (.A(_2624_),
    .B(_2643_),
    .C(_2644_),
    .Y(_2645_));
 sky130_fd_sc_hd__o21a_1 _7054_ (.A1(_2643_),
    .A2(_2644_),
    .B1(_2624_),
    .X(_2646_));
 sky130_fd_sc_hd__a211oi_2 _7055_ (.A1(_2436_),
    .A2(_2438_),
    .B1(_2645_),
    .C1(_2646_),
    .Y(_2647_));
 sky130_fd_sc_hd__o211a_1 _7056_ (.A1(_2645_),
    .A2(_2646_),
    .B1(_2436_),
    .C1(_2438_),
    .X(_2648_));
 sky130_fd_sc_hd__a211o_1 _7057_ (.A1(_2612_),
    .A2(_2613_),
    .B1(_2647_),
    .C1(_2648_),
    .X(_2649_));
 sky130_fd_sc_hd__o211ai_2 _7058_ (.A1(_2647_),
    .A2(_2648_),
    .B1(_2612_),
    .C1(_2613_),
    .Y(_2650_));
 sky130_fd_sc_hd__nand4_2 _7059_ (.A(_2610_),
    .B(_2611_),
    .C(_2649_),
    .D(_2650_),
    .Y(_2651_));
 sky130_fd_sc_hd__a22o_1 _7060_ (.A1(_2610_),
    .A2(_2611_),
    .B1(_2649_),
    .B2(_2650_),
    .X(_2652_));
 sky130_fd_sc_hd__o211a_1 _7061_ (.A1(_2502_),
    .A2(_2481_),
    .B1(_2651_),
    .C1(_2652_),
    .X(_2654_));
 sky130_fd_sc_hd__a211oi_1 _7062_ (.A1(_2651_),
    .A2(_2652_),
    .B1(_2502_),
    .C1(_2481_),
    .Y(_2655_));
 sky130_fd_sc_hd__nand2_1 _7063_ (.A(_2475_),
    .B(_2479_),
    .Y(_2656_));
 sky130_fd_sc_hd__nor3b_1 _7064_ (.A(_2654_),
    .B(_2655_),
    .C_N(_2656_),
    .Y(_2657_));
 sky130_fd_sc_hd__o21ba_1 _7065_ (.A1(_2654_),
    .A2(_2655_),
    .B1_N(_2656_),
    .X(_2658_));
 sky130_fd_sc_hd__or2_1 _7066_ (.A(_2657_),
    .B(_2658_),
    .X(_2659_));
 sky130_fd_sc_hd__a21oi_2 _7067_ (.A1(_2483_),
    .A2(_2485_),
    .B1(_2659_),
    .Y(_2660_));
 sky130_fd_sc_hd__and3_1 _7068_ (.A(_2483_),
    .B(_2485_),
    .C(_2659_),
    .X(_2661_));
 sky130_fd_sc_hd__nor2_1 _7069_ (.A(_2660_),
    .B(_2661_),
    .Y(_2662_));
 sky130_fd_sc_hd__nor2_1 _7070_ (.A(_2501_),
    .B(_2662_),
    .Y(_2663_));
 sky130_fd_sc_hd__and2_1 _7071_ (.A(_2501_),
    .B(_2662_),
    .X(_2665_));
 sky130_fd_sc_hd__or2_1 _7072_ (.A(_2663_),
    .B(_2665_),
    .X(_2666_));
 sky130_fd_sc_hd__a21oi_1 _7073_ (.A1(_2500_),
    .A2(_2497_),
    .B1(_2666_),
    .Y(_2667_));
 sky130_fd_sc_hd__a31o_1 _7074_ (.A1(_2500_),
    .A2(_2497_),
    .A3(_2666_),
    .B1(_3192_),
    .X(_2668_));
 sky130_fd_sc_hd__nor2_1 _7075_ (.A(_2667_),
    .B(_2668_),
    .Y(_2669_));
 sky130_fd_sc_hd__and2_2 _7076_ (.A(_2018_),
    .B(net54),
    .X(_2670_));
 sky130_fd_sc_hd__nor2_1 _7077_ (.A(_2018_),
    .B(net54),
    .Y(_2671_));
 sky130_fd_sc_hd__nor2_2 _7078_ (.A(_2670_),
    .B(_2671_),
    .Y(_2672_));
 sky130_fd_sc_hd__a21o_1 _7079_ (.A1(_2301_),
    .A2(_2306_),
    .B1(_2300_),
    .X(_2673_));
 sky130_fd_sc_hd__a21oi_1 _7080_ (.A1(_2672_),
    .A2(_2673_),
    .B1(_3596_),
    .Y(_2674_));
 sky130_fd_sc_hd__o21a_1 _7081_ (.A1(_2672_),
    .A2(_2673_),
    .B1(_2674_),
    .X(_2676_));
 sky130_fd_sc_hd__or2b_1 _7082_ (.A(_2299_),
    .B_N(_2007_),
    .X(_2677_));
 sky130_fd_sc_hd__a21o_1 _7083_ (.A1(_2311_),
    .A2(_2677_),
    .B1(_2672_),
    .X(_2678_));
 sky130_fd_sc_hd__a31oi_1 _7084_ (.A1(_2311_),
    .A2(_2672_),
    .A3(_2677_),
    .B1(_0181_),
    .Y(_2679_));
 sky130_fd_sc_hd__nor2_1 _7085_ (.A(_3589_),
    .B(_2670_),
    .Y(_2680_));
 sky130_fd_sc_hd__or2_1 _7086_ (.A(_2018_),
    .B(net54),
    .X(_2681_));
 sky130_fd_sc_hd__o21a_1 _7087_ (.A1(_1277_),
    .A2(_2680_),
    .B1(_2681_),
    .X(_2682_));
 sky130_fd_sc_hd__nor2_1 _7088_ (.A(_0848_),
    .B(_0196_),
    .Y(_2683_));
 sky130_fd_sc_hd__and2b_1 _7089_ (.A_N(_2683_),
    .B(_3161_),
    .X(_2684_));
 sky130_fd_sc_hd__a221o_1 _7090_ (.A1(_0854_),
    .A2(_2670_),
    .B1(_2671_),
    .B2(_0855_),
    .C1(_2684_),
    .X(_2685_));
 sky130_fd_sc_hd__mux4_1 _7091_ (.A0(_2018_),
    .A1(_2007_),
    .A2(_1821_),
    .A3(_1810_),
    .S0(_0863_),
    .S1(_0864_),
    .X(_2687_));
 sky130_fd_sc_hd__mux2_1 _7092_ (.A0(_1939_),
    .A1(_2687_),
    .S(_0866_),
    .X(_2688_));
 sky130_fd_sc_hd__mux4_1 _7093_ (.A0(_3097_),
    .A1(_0188_),
    .A2(_1284_),
    .A3(_2688_),
    .S0(_0867_),
    .S1(_0573_),
    .X(_2689_));
 sky130_fd_sc_hd__a2bb2o_1 _7094_ (.A1_N(_3156_),
    .A2_N(_0201_),
    .B1(_2689_),
    .B2(_0844_),
    .X(_2690_));
 sky130_fd_sc_hd__or3_1 _7095_ (.A(_2682_),
    .B(_2685_),
    .C(_2690_),
    .X(_2691_));
 sky130_fd_sc_hd__a21oi_1 _7096_ (.A1(_2678_),
    .A2(_2679_),
    .B1(_2691_),
    .Y(_2692_));
 sky130_fd_sc_hd__or3b_1 _7097_ (.A(_2669_),
    .B(_2676_),
    .C_N(_2692_),
    .X(_2693_));
 sky130_fd_sc_hd__clkbuf_1 _7098_ (.A(_2693_),
    .X(net90));
 sky130_fd_sc_hd__nor2_1 _7099_ (.A(_2051_),
    .B(net56),
    .Y(_2694_));
 sky130_fd_sc_hd__and2_1 _7100_ (.A(_2051_),
    .B(net56),
    .X(_2695_));
 sky130_fd_sc_hd__nor2_2 _7101_ (.A(_2694_),
    .B(_2695_),
    .Y(_2697_));
 sky130_fd_sc_hd__and2_1 _7102_ (.A(_2681_),
    .B(_2673_),
    .X(_2698_));
 sky130_fd_sc_hd__or3_1 _7103_ (.A(_2670_),
    .B(_2697_),
    .C(_2698_),
    .X(_2699_));
 sky130_fd_sc_hd__o21ai_2 _7104_ (.A1(_2670_),
    .A2(_2698_),
    .B1(_2697_),
    .Y(_2700_));
 sky130_fd_sc_hd__or2b_1 _7105_ (.A(net54),
    .B_N(_2018_),
    .X(_2701_));
 sky130_fd_sc_hd__nand3_1 _7106_ (.A(_2678_),
    .B(_2697_),
    .C(_2701_),
    .Y(_2702_));
 sky130_fd_sc_hd__a21o_1 _7107_ (.A1(_2678_),
    .A2(_2701_),
    .B1(_2697_),
    .X(_2703_));
 sky130_fd_sc_hd__and4bb_1 _7108_ (.A_N(_2564_),
    .B_N(_2566_),
    .C(_2605_),
    .D(_2606_),
    .X(_2704_));
 sky130_fd_sc_hd__o211a_1 _7109_ (.A1(_2353_),
    .A2(_2503_),
    .B1(_2534_),
    .C1(_2535_),
    .X(_2705_));
 sky130_fd_sc_hd__and4_1 _7110_ (.A(_2536_),
    .B(_2537_),
    .C(_2560_),
    .D(_2561_),
    .X(_2706_));
 sky130_fd_sc_hd__nor3_2 _7111_ (.A(_2522_),
    .B(_2523_),
    .C(_2533_),
    .Y(_2708_));
 sky130_fd_sc_hd__a22o_1 _7112_ (.A1(_0521_),
    .A2(net22),
    .B1(net24),
    .B2(_0881_),
    .X(_2709_));
 sky130_fd_sc_hd__nand4_2 _7113_ (.A(_0881_),
    .B(_0521_),
    .C(net22),
    .D(_2051_),
    .Y(_2710_));
 sky130_fd_sc_hd__a22o_1 _7114_ (.A1(_0980_),
    .A2(net21),
    .B1(_2709_),
    .B2(_2710_),
    .X(_2711_));
 sky130_fd_sc_hd__nand4_2 _7115_ (.A(_0980_),
    .B(net21),
    .C(_2709_),
    .D(_2710_),
    .Y(_2712_));
 sky130_fd_sc_hd__a21bo_1 _7116_ (.A1(_2504_),
    .A2(_2506_),
    .B1_N(_2505_),
    .X(_2713_));
 sky130_fd_sc_hd__nand3_1 _7117_ (.A(_2711_),
    .B(_2712_),
    .C(_2713_),
    .Y(_2714_));
 sky130_fd_sc_hd__a21o_1 _7118_ (.A1(_2711_),
    .A2(_2712_),
    .B1(_2713_),
    .X(_2715_));
 sky130_fd_sc_hd__a22oi_1 _7119_ (.A1(_0063_),
    .A2(_1799_),
    .B1(net20),
    .B2(_0183_),
    .Y(_2716_));
 sky130_fd_sc_hd__and4_1 _7120_ (.A(_0172_),
    .B(_0052_),
    .C(_1799_),
    .D(net20),
    .X(_2717_));
 sky130_fd_sc_hd__nor2_1 _7121_ (.A(_2716_),
    .B(_2717_),
    .Y(_2719_));
 sky130_fd_sc_hd__nand2_1 _7122_ (.A(_2903_),
    .B(_1767_),
    .Y(_2720_));
 sky130_fd_sc_hd__xnor2_1 _7123_ (.A(_2719_),
    .B(_2720_),
    .Y(_2721_));
 sky130_fd_sc_hd__nand3_1 _7124_ (.A(_2714_),
    .B(_2715_),
    .C(_2721_),
    .Y(_2722_));
 sky130_fd_sc_hd__a21o_1 _7125_ (.A1(_2714_),
    .A2(_2715_),
    .B1(_2721_),
    .X(_2723_));
 sky130_fd_sc_hd__a21bo_1 _7126_ (.A1(_2512_),
    .A2(_2517_),
    .B1_N(_2511_),
    .X(_2724_));
 sky130_fd_sc_hd__and3_1 _7127_ (.A(_2722_),
    .B(_2723_),
    .C(_2724_),
    .X(_2725_));
 sky130_fd_sc_hd__a21oi_1 _7128_ (.A1(_2722_),
    .A2(_2723_),
    .B1(_2724_),
    .Y(_2726_));
 sky130_fd_sc_hd__a31o_1 _7129_ (.A1(_3386_),
    .A2(_1898_),
    .A3(_2528_),
    .B1(_2527_),
    .X(_2727_));
 sky130_fd_sc_hd__a31o_1 _7130_ (.A1(_2903_),
    .A2(_1745_),
    .A3(_2515_),
    .B1(_2514_),
    .X(_2728_));
 sky130_fd_sc_hd__nand2_1 _7131_ (.A(_3386_),
    .B(_1931_),
    .Y(_2730_));
 sky130_fd_sc_hd__a22oi_1 _7132_ (.A1(_3273_),
    .A2(_1952_),
    .B1(_1745_),
    .B2(_3198_),
    .Y(_2731_));
 sky130_fd_sc_hd__and4_1 _7133_ (.A(_3198_),
    .B(_3273_),
    .C(_1952_),
    .D(_1745_),
    .X(_2732_));
 sky130_fd_sc_hd__nor2_1 _7134_ (.A(_2731_),
    .B(_2732_),
    .Y(_2733_));
 sky130_fd_sc_hd__xnor2_1 _7135_ (.A(_2730_),
    .B(_2733_),
    .Y(_2734_));
 sky130_fd_sc_hd__xor2_1 _7136_ (.A(_2728_),
    .B(_2734_),
    .X(_2735_));
 sky130_fd_sc_hd__xnor2_1 _7137_ (.A(_2727_),
    .B(_2735_),
    .Y(_2736_));
 sky130_fd_sc_hd__or3_2 _7138_ (.A(_2725_),
    .B(_2726_),
    .C(_2736_),
    .X(_2737_));
 sky130_fd_sc_hd__o21ai_2 _7139_ (.A1(_2725_),
    .A2(_2726_),
    .B1(_2736_),
    .Y(_2738_));
 sky130_fd_sc_hd__o211ai_4 _7140_ (.A1(_2522_),
    .A2(_2708_),
    .B1(_2737_),
    .C1(_2738_),
    .Y(_2739_));
 sky130_fd_sc_hd__a211o_1 _7141_ (.A1(_2737_),
    .A2(_2738_),
    .B1(_2522_),
    .C1(_2708_),
    .X(_2741_));
 sky130_fd_sc_hd__and2_1 _7142_ (.A(_2525_),
    .B(_2530_),
    .X(_2742_));
 sky130_fd_sc_hd__and2_1 _7143_ (.A(_2524_),
    .B(_2531_),
    .X(_2743_));
 sky130_fd_sc_hd__a22oi_2 _7144_ (.A1(_0174_),
    .A2(_2543_),
    .B1(_2576_),
    .B2(_3720_),
    .Y(_2744_));
 sky130_fd_sc_hd__and4_1 _7145_ (.A(_3720_),
    .B(_0174_),
    .C(_2543_),
    .D(_2576_),
    .X(_2745_));
 sky130_fd_sc_hd__or2_1 _7146_ (.A(_2744_),
    .B(_2745_),
    .X(_2746_));
 sky130_fd_sc_hd__nand2_1 _7147_ (.A(_0293_),
    .B(_2510_),
    .Y(_2747_));
 sky130_fd_sc_hd__xnor2_1 _7148_ (.A(_2746_),
    .B(_2747_),
    .Y(_2748_));
 sky130_fd_sc_hd__a22oi_1 _7149_ (.A1(_3513_),
    .A2(_1865_),
    .B1(_1898_),
    .B2(_3425_),
    .Y(_2749_));
 sky130_fd_sc_hd__and4_1 _7150_ (.A(_3425_),
    .B(_3513_),
    .C(_1865_),
    .D(_1898_),
    .X(_2750_));
 sky130_fd_sc_hd__nor2_1 _7151_ (.A(_2749_),
    .B(_2750_),
    .Y(_2752_));
 sky130_fd_sc_hd__nand2_1 _7152_ (.A(_3685_),
    .B(_2609_),
    .Y(_2753_));
 sky130_fd_sc_hd__xnor2_1 _7153_ (.A(_2752_),
    .B(_2753_),
    .Y(_2754_));
 sky130_fd_sc_hd__nand2_1 _7154_ (.A(_2549_),
    .B(_2551_),
    .Y(_2755_));
 sky130_fd_sc_hd__xnor2_1 _7155_ (.A(_2754_),
    .B(_2755_),
    .Y(_2756_));
 sky130_fd_sc_hd__xor2_1 _7156_ (.A(_2748_),
    .B(_2756_),
    .X(_2757_));
 sky130_fd_sc_hd__o21a_2 _7157_ (.A1(_2742_),
    .A2(_2743_),
    .B1(_2757_),
    .X(_2758_));
 sky130_fd_sc_hd__nor3_2 _7158_ (.A(_2742_),
    .B(_2743_),
    .C(_2757_),
    .Y(_2759_));
 sky130_fd_sc_hd__a211o_1 _7159_ (.A1(_2553_),
    .A2(_2556_),
    .B1(_2758_),
    .C1(_2759_),
    .X(_2760_));
 sky130_fd_sc_hd__o211ai_4 _7160_ (.A1(_2758_),
    .A2(_2759_),
    .B1(_2553_),
    .C1(_2556_),
    .Y(_2761_));
 sky130_fd_sc_hd__nand4_4 _7161_ (.A(_2739_),
    .B(_2741_),
    .C(_2760_),
    .D(_2761_),
    .Y(_2763_));
 sky130_fd_sc_hd__a22o_1 _7162_ (.A1(_2739_),
    .A2(_2741_),
    .B1(_2760_),
    .B2(_2761_),
    .X(_2764_));
 sky130_fd_sc_hd__o211ai_4 _7163_ (.A1(_2705_),
    .A2(_2706_),
    .B1(_2763_),
    .C1(_2764_),
    .Y(_2765_));
 sky130_fd_sc_hd__a211o_1 _7164_ (.A1(_2763_),
    .A2(_2764_),
    .B1(_2705_),
    .C1(_2706_),
    .X(_2766_));
 sky130_fd_sc_hd__a21bo_1 _7165_ (.A1(_2586_),
    .A2(_2600_),
    .B1_N(_2599_),
    .X(_2767_));
 sky130_fd_sc_hd__and2b_1 _7166_ (.A_N(_2558_),
    .B(_2560_),
    .X(_2768_));
 sky130_fd_sc_hd__a22oi_1 _7167_ (.A1(_2171_),
    .A2(_1170_),
    .B1(_1295_),
    .B2(_2127_),
    .Y(_2769_));
 sky130_fd_sc_hd__and4_1 _7168_ (.A(_2127_),
    .B(_2171_),
    .C(_1170_),
    .D(_1295_),
    .X(_2770_));
 sky130_fd_sc_hd__nor2_1 _7169_ (.A(_2769_),
    .B(_2770_),
    .Y(_2771_));
 sky130_fd_sc_hd__nand2_1 _7170_ (.A(_2456_),
    .B(_1448_),
    .Y(_2772_));
 sky130_fd_sc_hd__xor2_1 _7171_ (.A(_2771_),
    .B(_2772_),
    .X(_2774_));
 sky130_fd_sc_hd__a22o_1 _7172_ (.A1(_2664_),
    .A2(_0722_),
    .B1(_0875_),
    .B2(_2270_),
    .X(_2775_));
 sky130_fd_sc_hd__nand4_1 _7173_ (.A(_2270_),
    .B(_2664_),
    .C(_0722_),
    .D(_0875_),
    .Y(_2776_));
 sky130_fd_sc_hd__nand2_1 _7174_ (.A(_2775_),
    .B(_2776_),
    .Y(_2777_));
 sky130_fd_sc_hd__nand2_1 _7175_ (.A(_2226_),
    .B(_1008_),
    .Y(_2778_));
 sky130_fd_sc_hd__xor2_1 _7176_ (.A(_2777_),
    .B(_2778_),
    .X(_2779_));
 sky130_fd_sc_hd__or2_1 _7177_ (.A(_2578_),
    .B(_2580_),
    .X(_2780_));
 sky130_fd_sc_hd__xnor2_1 _7178_ (.A(_2779_),
    .B(_2780_),
    .Y(_2781_));
 sky130_fd_sc_hd__nor2_1 _7179_ (.A(_2774_),
    .B(_2781_),
    .Y(_2782_));
 sky130_fd_sc_hd__and2_1 _7180_ (.A(_2774_),
    .B(_2781_),
    .X(_2783_));
 sky130_fd_sc_hd__nor2_1 _7181_ (.A(_2782_),
    .B(_2783_),
    .Y(_2785_));
 sky130_fd_sc_hd__nand2_1 _7182_ (.A(_2591_),
    .B(_2593_),
    .Y(_2786_));
 sky130_fd_sc_hd__o2bb2a_1 _7183_ (.A1_N(_2543_),
    .A2_N(_2542_),
    .B1(_2545_),
    .B2(_2546_),
    .X(_2787_));
 sky130_fd_sc_hd__nand2_1 _7184_ (.A(_2762_),
    .B(_0454_),
    .Y(_2788_));
 sky130_fd_sc_hd__xnor2_1 _7185_ (.A(_0420_),
    .B(_2788_),
    .Y(_2789_));
 sky130_fd_sc_hd__nand2_1 _7186_ (.A(_2718_),
    .B(_0689_),
    .Y(_2790_));
 sky130_fd_sc_hd__xor2_1 _7187_ (.A(_2789_),
    .B(_2790_),
    .X(_2791_));
 sky130_fd_sc_hd__xor2_1 _7188_ (.A(_2787_),
    .B(_2791_),
    .X(_2792_));
 sky130_fd_sc_hd__xnor2_1 _7189_ (.A(_2786_),
    .B(_2792_),
    .Y(_2793_));
 sky130_fd_sc_hd__a21bo_1 _7190_ (.A1(_2589_),
    .A2(_2595_),
    .B1_N(_2594_),
    .X(_2794_));
 sky130_fd_sc_hd__xnor2_1 _7191_ (.A(_2793_),
    .B(_2794_),
    .Y(_2796_));
 sky130_fd_sc_hd__xnor2_1 _7192_ (.A(_2785_),
    .B(_2796_),
    .Y(_2797_));
 sky130_fd_sc_hd__xor2_1 _7193_ (.A(_2768_),
    .B(_2797_),
    .X(_2798_));
 sky130_fd_sc_hd__xor2_1 _7194_ (.A(_2767_),
    .B(_2798_),
    .X(_2799_));
 sky130_fd_sc_hd__nand3_1 _7195_ (.A(_2765_),
    .B(_2766_),
    .C(_2799_),
    .Y(_2800_));
 sky130_fd_sc_hd__a21o_1 _7196_ (.A1(_2765_),
    .A2(_2766_),
    .B1(_2799_),
    .X(_2801_));
 sky130_fd_sc_hd__o211a_1 _7197_ (.A1(_2564_),
    .A2(_2704_),
    .B1(_2800_),
    .C1(_2801_),
    .X(_2802_));
 sky130_fd_sc_hd__a211oi_2 _7198_ (.A1(_2800_),
    .A2(_2801_),
    .B1(_2564_),
    .C1(_2704_),
    .Y(_2803_));
 sky130_fd_sc_hd__inv_2 _7199_ (.A(_2643_),
    .Y(_2804_));
 sky130_fd_sc_hd__or3_1 _7200_ (.A(_2624_),
    .B(_2643_),
    .C(_2644_),
    .X(_2805_));
 sky130_fd_sc_hd__a22oi_1 _7201_ (.A1(_0226_),
    .A2(_2263_),
    .B1(_2299_),
    .B2(_1045_),
    .Y(_2807_));
 sky130_fd_sc_hd__and4_1 _7202_ (.A(_0226_),
    .B(_1045_),
    .C(net52),
    .D(_2299_),
    .X(_2808_));
 sky130_fd_sc_hd__nor2_1 _7203_ (.A(_2807_),
    .B(_2808_),
    .Y(_2809_));
 sky130_fd_sc_hd__nand2_1 _7204_ (.A(_1056_),
    .B(net54),
    .Y(_2810_));
 sky130_fd_sc_hd__xor2_1 _7205_ (.A(_2809_),
    .B(_2810_),
    .X(_2811_));
 sky130_fd_sc_hd__or2_1 _7206_ (.A(_2617_),
    .B(_2619_),
    .X(_2812_));
 sky130_fd_sc_hd__and2b_1 _7207_ (.A_N(_2811_),
    .B(_2812_),
    .X(_2813_));
 sky130_fd_sc_hd__and2b_1 _7208_ (.A_N(_2812_),
    .B(_2811_),
    .X(_2814_));
 sky130_fd_sc_hd__or2_1 _7209_ (.A(_2813_),
    .B(_2814_),
    .X(_2815_));
 sky130_fd_sc_hd__nand2_1 _7210_ (.A(_3209_),
    .B(net56),
    .Y(_2816_));
 sky130_fd_sc_hd__xor2_1 _7211_ (.A(_2815_),
    .B(_2816_),
    .X(_2818_));
 sky130_fd_sc_hd__nand2_1 _7212_ (.A(_2622_),
    .B(_2818_),
    .Y(_2819_));
 sky130_fd_sc_hd__or2_1 _7213_ (.A(_2622_),
    .B(_2818_),
    .X(_2820_));
 sky130_fd_sc_hd__nand2_1 _7214_ (.A(_2819_),
    .B(_2820_),
    .Y(_2821_));
 sky130_fd_sc_hd__or2b_1 _7215_ (.A(_2635_),
    .B_N(_2629_),
    .X(_2822_));
 sky130_fd_sc_hd__nand2_1 _7216_ (.A(_2628_),
    .B(_2636_),
    .Y(_2823_));
 sky130_fd_sc_hd__nand2_1 _7217_ (.A(_2581_),
    .B(_2582_),
    .Y(_2824_));
 sky130_fd_sc_hd__a41o_1 _7218_ (.A1(_1023_),
    .A2(_2346_),
    .A3(_1608_),
    .A4(_1797_),
    .B1(_2634_),
    .X(_2825_));
 sky130_fd_sc_hd__or2_1 _7219_ (.A(_2572_),
    .B(_2574_),
    .X(_2826_));
 sky130_fd_sc_hd__a22oi_1 _7220_ (.A1(_2401_),
    .A2(_1608_),
    .B1(_1797_),
    .B2(_2335_),
    .Y(_2827_));
 sky130_fd_sc_hd__and4_1 _7221_ (.A(_2335_),
    .B(_2401_),
    .C(_1607_),
    .D(_1797_),
    .X(_2829_));
 sky130_fd_sc_hd__nand2_1 _7222_ (.A(_0117_),
    .B(_1949_),
    .Y(_2830_));
 sky130_fd_sc_hd__o21ai_1 _7223_ (.A1(_2827_),
    .A2(_2829_),
    .B1(_2830_),
    .Y(_2831_));
 sky130_fd_sc_hd__or3_1 _7224_ (.A(_2827_),
    .B(_2829_),
    .C(_2830_),
    .X(_2832_));
 sky130_fd_sc_hd__nand2_1 _7225_ (.A(_2831_),
    .B(_2832_),
    .Y(_2833_));
 sky130_fd_sc_hd__xnor2_1 _7226_ (.A(_2826_),
    .B(_2833_),
    .Y(_2834_));
 sky130_fd_sc_hd__xnor2_1 _7227_ (.A(_2825_),
    .B(_2834_),
    .Y(_2835_));
 sky130_fd_sc_hd__a21oi_2 _7228_ (.A1(_2824_),
    .A2(_2584_),
    .B1(_2835_),
    .Y(_2836_));
 sky130_fd_sc_hd__and3_1 _7229_ (.A(_2824_),
    .B(_2584_),
    .C(_2835_),
    .X(_2837_));
 sky130_fd_sc_hd__a211o_1 _7230_ (.A1(_2822_),
    .A2(_2823_),
    .B1(_2836_),
    .C1(_2837_),
    .X(_2838_));
 sky130_fd_sc_hd__o211ai_2 _7231_ (.A1(_2836_),
    .A2(_2837_),
    .B1(_2822_),
    .C1(_2823_),
    .Y(_2840_));
 sky130_fd_sc_hd__o211a_1 _7232_ (.A1(_2638_),
    .A2(_2640_),
    .B1(_2838_),
    .C1(_2840_),
    .X(_2841_));
 sky130_fd_sc_hd__a211oi_2 _7233_ (.A1(_2838_),
    .A2(_2840_),
    .B1(_2638_),
    .C1(_2640_),
    .Y(_2842_));
 sky130_fd_sc_hd__nor3_2 _7234_ (.A(_2821_),
    .B(_2841_),
    .C(_2842_),
    .Y(_2843_));
 sky130_fd_sc_hd__o21a_1 _7235_ (.A1(_2841_),
    .A2(_2842_),
    .B1(_2821_),
    .X(_2844_));
 sky130_fd_sc_hd__a211oi_4 _7236_ (.A1(_2603_),
    .A2(_2605_),
    .B1(_2843_),
    .C1(_2844_),
    .Y(_2845_));
 sky130_fd_sc_hd__o211a_1 _7237_ (.A1(_2843_),
    .A2(_2844_),
    .B1(_2603_),
    .C1(_2605_),
    .X(_2846_));
 sky130_fd_sc_hd__a211oi_2 _7238_ (.A1(_2804_),
    .A2(_2805_),
    .B1(_2845_),
    .C1(_2846_),
    .Y(_2847_));
 sky130_fd_sc_hd__o211a_1 _7239_ (.A1(_2845_),
    .A2(_2846_),
    .B1(_2804_),
    .C1(_2805_),
    .X(_2848_));
 sky130_fd_sc_hd__nor4_1 _7240_ (.A(_2802_),
    .B(_2803_),
    .C(_2847_),
    .D(_2848_),
    .Y(_2849_));
 sky130_fd_sc_hd__o22a_1 _7241_ (.A1(_2802_),
    .A2(_2803_),
    .B1(_2847_),
    .B2(_2848_),
    .X(_2851_));
 sky130_fd_sc_hd__a211oi_1 _7242_ (.A1(_2610_),
    .A2(_2651_),
    .B1(net197),
    .C1(_2851_),
    .Y(_2852_));
 sky130_fd_sc_hd__o211ai_1 _7243_ (.A1(net197),
    .A2(_2851_),
    .B1(_2610_),
    .C1(_2651_),
    .Y(_2853_));
 sky130_fd_sc_hd__and2b_1 _7244_ (.A_N(_2852_),
    .B(_2853_),
    .X(_2854_));
 sky130_fd_sc_hd__or2b_1 _7245_ (.A(_2647_),
    .B_N(_2649_),
    .X(_2855_));
 sky130_fd_sc_hd__xor2_1 _7246_ (.A(_2854_),
    .B(_2855_),
    .X(_2856_));
 sky130_fd_sc_hd__o21ai_1 _7247_ (.A1(_2654_),
    .A2(_2657_),
    .B1(_2856_),
    .Y(_2857_));
 sky130_fd_sc_hd__or3_1 _7248_ (.A(_2654_),
    .B(_2657_),
    .C(_2856_),
    .X(_2858_));
 sky130_fd_sc_hd__and2_1 _7249_ (.A(_2857_),
    .B(_2858_),
    .X(_2859_));
 sky130_fd_sc_hd__nand2_1 _7250_ (.A(_2660_),
    .B(_2859_),
    .Y(_2860_));
 sky130_fd_sc_hd__or2_1 _7251_ (.A(_2660_),
    .B(_2859_),
    .X(_2862_));
 sky130_fd_sc_hd__nand2_1 _7252_ (.A(_2860_),
    .B(_2862_),
    .Y(_2863_));
 sky130_fd_sc_hd__nand2_1 _7253_ (.A(_2487_),
    .B(_2500_),
    .Y(_2864_));
 sky130_fd_sc_hd__o2bb2a_1 _7254_ (.A1_N(_2864_),
    .A2_N(_2662_),
    .B1(_2497_),
    .B2(_2663_),
    .X(_2865_));
 sky130_fd_sc_hd__o21ai_1 _7255_ (.A1(_2863_),
    .A2(_2865_),
    .B1(_0320_),
    .Y(_2866_));
 sky130_fd_sc_hd__a21oi_1 _7256_ (.A1(_2863_),
    .A2(_2865_),
    .B1(_2866_),
    .Y(_2867_));
 sky130_fd_sc_hd__mux4_1 _7257_ (.A0(_2051_),
    .A1(_2018_),
    .A2(_2007_),
    .A3(_1821_),
    .S0(_0863_),
    .S1(_0864_),
    .X(_2868_));
 sky130_fd_sc_hd__mux2_1 _7258_ (.A0(_2114_),
    .A1(_2868_),
    .S(_0866_),
    .X(_2869_));
 sky130_fd_sc_hd__mux4_1 _7259_ (.A0(_3213_),
    .A1(_0305_),
    .A2(_1309_),
    .A3(_2869_),
    .S0(_0867_),
    .S1(_0573_),
    .X(_2870_));
 sky130_fd_sc_hd__nand2_1 _7260_ (.A(_2051_),
    .B(net56),
    .Y(_2871_));
 sky130_fd_sc_hd__a21oi_1 _7261_ (.A1(_0438_),
    .A2(_2871_),
    .B1(_1277_),
    .Y(_2872_));
 sky130_fd_sc_hd__nor2_1 _7262_ (.A(_2694_),
    .B(_2872_),
    .Y(_2873_));
 sky130_fd_sc_hd__mux2_1 _7263_ (.A0(_0571_),
    .A1(_2062_),
    .S(_2683_),
    .X(_2874_));
 sky130_fd_sc_hd__nor2_1 _7264_ (.A(_0313_),
    .B(_2319_),
    .Y(_2875_));
 sky130_fd_sc_hd__a22o_1 _7265_ (.A1(_0855_),
    .A2(_2694_),
    .B1(_2695_),
    .B2(_0854_),
    .X(_2876_));
 sky130_fd_sc_hd__a211o_1 _7266_ (.A1(_0575_),
    .A2(_2874_),
    .B1(_2875_),
    .C1(_2876_),
    .X(_2877_));
 sky130_fd_sc_hd__a211o_1 _7267_ (.A1(_0844_),
    .A2(_2870_),
    .B1(_2873_),
    .C1(_2877_),
    .X(_2878_));
 sky130_fd_sc_hd__a311o_1 _7268_ (.A1(_3571_),
    .A2(_2702_),
    .A3(_2703_),
    .B1(_2867_),
    .C1(_2878_),
    .X(_2879_));
 sky130_fd_sc_hd__a31o_4 _7269_ (.A1(_0419_),
    .A2(_2699_),
    .A3(_2700_),
    .B1(_2879_),
    .X(net92));
 sky130_fd_sc_hd__or2_1 _7270_ (.A(_0571_),
    .B(net57),
    .X(_2880_));
 sky130_fd_sc_hd__nand2_1 _7271_ (.A(_0571_),
    .B(net57),
    .Y(_2882_));
 sky130_fd_sc_hd__nand2_2 _7272_ (.A(_2880_),
    .B(_2882_),
    .Y(_2883_));
 sky130_fd_sc_hd__a21oi_1 _7273_ (.A1(_2871_),
    .A2(_2700_),
    .B1(_2883_),
    .Y(_2884_));
 sky130_fd_sc_hd__a31o_1 _7274_ (.A1(_2871_),
    .A2(_2700_),
    .A3(_2883_),
    .B1(_3596_),
    .X(_2885_));
 sky130_fd_sc_hd__or2_1 _7275_ (.A(_2884_),
    .B(_2885_),
    .X(_2886_));
 sky130_fd_sc_hd__or2b_1 _7276_ (.A(net56),
    .B_N(_2051_),
    .X(_2887_));
 sky130_fd_sc_hd__and3b_1 _7277_ (.A_N(_2883_),
    .B(_2887_),
    .C(_2703_),
    .X(_2888_));
 sky130_fd_sc_hd__a21boi_1 _7278_ (.A1(_2703_),
    .A2(_2887_),
    .B1_N(_2883_),
    .Y(_2889_));
 sky130_fd_sc_hd__mux4_1 _7279_ (.A0(_0571_),
    .A1(_2018_),
    .A2(_2051_),
    .A3(_2007_),
    .S0(_0864_),
    .S1(_0863_),
    .X(_2890_));
 sky130_fd_sc_hd__mux2_1 _7280_ (.A0(_2285_),
    .A1(_2890_),
    .S(_0866_),
    .X(_2891_));
 sky130_fd_sc_hd__mux4_1 _7281_ (.A0(_3285_),
    .A1(_0435_),
    .A2(_1467_),
    .A3(_2891_),
    .S0(_0867_),
    .S1(_0573_),
    .X(_2893_));
 sky130_fd_sc_hd__nand2_1 _7282_ (.A(_0844_),
    .B(_2893_),
    .Y(_2894_));
 sky130_fd_sc_hd__o22a_1 _7283_ (.A1(_0309_),
    .A2(_2882_),
    .B1(_2883_),
    .B2(_3589_),
    .X(_2895_));
 sky130_fd_sc_hd__nand2_1 _7284_ (.A(_1277_),
    .B(_2880_),
    .Y(_2896_));
 sky130_fd_sc_hd__o21ba_1 _7285_ (.A1(_3712_),
    .A2(_2880_),
    .B1_N(_3161_),
    .X(_2897_));
 sky130_fd_sc_hd__and3_1 _7286_ (.A(_2895_),
    .B(_2896_),
    .C(_2897_),
    .X(_2898_));
 sky130_fd_sc_hd__o311a_1 _7287_ (.A1(_3144_),
    .A2(_0196_),
    .A3(_2319_),
    .B1(_2894_),
    .C1(_2898_),
    .X(_2899_));
 sky130_fd_sc_hd__o21ai_1 _7288_ (.A1(_2863_),
    .A2(_2865_),
    .B1(_2860_),
    .Y(_2900_));
 sky130_fd_sc_hd__nand2_1 _7289_ (.A(_1067_),
    .B(net56),
    .Y(_2901_));
 sky130_fd_sc_hd__a31o_1 _7290_ (.A1(_3685_),
    .A2(_0862_),
    .A3(_2752_),
    .B1(_2750_),
    .X(_2902_));
 sky130_fd_sc_hd__nor2_1 _7291_ (.A(_2768_),
    .B(_2797_),
    .Y(_2904_));
 sky130_fd_sc_hd__a21o_1 _7292_ (.A1(_2767_),
    .A2(_2798_),
    .B1(_2904_),
    .X(_2905_));
 sky130_fd_sc_hd__xor2_1 _7293_ (.A(_2902_),
    .B(_2905_),
    .X(_2906_));
 sky130_fd_sc_hd__xor2_1 _7294_ (.A(_2901_),
    .B(_2906_),
    .X(_2907_));
 sky130_fd_sc_hd__a211oi_2 _7295_ (.A1(_2553_),
    .A2(_2556_),
    .B1(_2758_),
    .C1(_2759_),
    .Y(_2908_));
 sky130_fd_sc_hd__a211oi_1 _7296_ (.A1(_3137_),
    .A2(_1008_),
    .B1(_2758_),
    .C1(_2908_),
    .Y(_2909_));
 sky130_fd_sc_hd__o211a_1 _7297_ (.A1(_2758_),
    .A2(_2908_),
    .B1(_3137_),
    .C1(_1008_),
    .X(_2910_));
 sky130_fd_sc_hd__nor2_1 _7298_ (.A(_2909_),
    .B(_2910_),
    .Y(_2911_));
 sky130_fd_sc_hd__xnor2_1 _7299_ (.A(_2907_),
    .B(_2911_),
    .Y(_2912_));
 sky130_fd_sc_hd__o211a_1 _7300_ (.A1(_2802_),
    .A2(net102),
    .B1(_3139_),
    .C1(_1608_),
    .X(_2913_));
 sky130_fd_sc_hd__a211oi_1 _7301_ (.A1(_3139_),
    .A2(_1608_),
    .B1(_2802_),
    .C1(net102),
    .Y(_2915_));
 sky130_fd_sc_hd__nor2_1 _7302_ (.A(_2913_),
    .B(_2915_),
    .Y(_2916_));
 sky130_fd_sc_hd__o211a_1 _7303_ (.A1(_2845_),
    .A2(_2847_),
    .B1(_1023_),
    .C1(_2263_),
    .X(_2917_));
 sky130_fd_sc_hd__a211oi_1 _7304_ (.A1(_1023_),
    .A2(_2263_),
    .B1(_2845_),
    .C1(_2847_),
    .Y(_2918_));
 sky130_fd_sc_hd__nor2_1 _7305_ (.A(_2917_),
    .B(_2918_),
    .Y(_2919_));
 sky130_fd_sc_hd__a211oi_1 _7306_ (.A1(_1034_),
    .A2(_2299_),
    .B1(_2841_),
    .C1(_2843_),
    .Y(_2920_));
 sky130_fd_sc_hd__o211a_1 _7307_ (.A1(_2841_),
    .A2(_2843_),
    .B1(_1034_),
    .C1(_2299_),
    .X(_2921_));
 sky130_fd_sc_hd__nor2_1 _7308_ (.A(_2920_),
    .B(_2921_),
    .Y(_2922_));
 sky130_fd_sc_hd__o21bai_2 _7309_ (.A1(_2744_),
    .A2(_2747_),
    .B1_N(_2745_),
    .Y(_2923_));
 sky130_fd_sc_hd__nand2_1 _7310_ (.A(_0328_),
    .B(_0558_),
    .Y(_2924_));
 sky130_fd_sc_hd__xnor2_2 _7311_ (.A(_2923_),
    .B(_2924_),
    .Y(_2926_));
 sky130_fd_sc_hd__xnor2_1 _7312_ (.A(_2922_),
    .B(_2926_),
    .Y(_2927_));
 sky130_fd_sc_hd__xnor2_1 _7313_ (.A(_2919_),
    .B(_2927_),
    .Y(_2928_));
 sky130_fd_sc_hd__xnor2_1 _7314_ (.A(_2916_),
    .B(_2928_),
    .Y(_2929_));
 sky130_fd_sc_hd__xnor2_1 _7315_ (.A(_2912_),
    .B(_2929_),
    .Y(_2930_));
 sky130_fd_sc_hd__a31o_1 _7316_ (.A1(_3139_),
    .A2(_1448_),
    .A3(_2771_),
    .B1(_2770_),
    .X(_2931_));
 sky130_fd_sc_hd__nand2_1 _7317_ (.A(_0174_),
    .B(_2587_),
    .Y(_2932_));
 sky130_fd_sc_hd__nand2_1 _7318_ (.A(_2675_),
    .B(_0875_),
    .Y(_2933_));
 sky130_fd_sc_hd__nand2_1 _7319_ (.A(_3133_),
    .B(_0722_),
    .Y(_2934_));
 sky130_fd_sc_hd__xor2_1 _7320_ (.A(_2933_),
    .B(_2934_),
    .X(_2935_));
 sky130_fd_sc_hd__xnor2_1 _7321_ (.A(_2932_),
    .B(_2935_),
    .Y(_2937_));
 sky130_fd_sc_hd__a32o_1 _7322_ (.A1(_2826_),
    .A2(_2831_),
    .A3(_2832_),
    .B1(_2834_),
    .B2(_2825_),
    .X(_2938_));
 sky130_fd_sc_hd__nand2_1 _7323_ (.A(_3198_),
    .B(_1778_),
    .Y(_2939_));
 sky130_fd_sc_hd__nand2_1 _7324_ (.A(_3685_),
    .B(_1876_),
    .Y(_2940_));
 sky130_fd_sc_hd__nand2_1 _7325_ (.A(_2714_),
    .B(_2722_),
    .Y(_2941_));
 sky130_fd_sc_hd__xor2_1 _7326_ (.A(_2940_),
    .B(_2941_),
    .X(_2942_));
 sky130_fd_sc_hd__xnor2_1 _7327_ (.A(_2939_),
    .B(_2942_),
    .Y(_2943_));
 sky130_fd_sc_hd__nand2_1 _7328_ (.A(_3273_),
    .B(_1756_),
    .Y(_2944_));
 sky130_fd_sc_hd__a21oi_1 _7329_ (.A1(_3198_),
    .A2(_1963_),
    .B1(_2944_),
    .Y(_2945_));
 sky130_fd_sc_hd__or3_1 _7330_ (.A(_2730_),
    .B(_2731_),
    .C(_2732_),
    .X(_2946_));
 sky130_fd_sc_hd__mux2_1 _7331_ (.A0(_2944_),
    .A1(_2945_),
    .S(_2946_),
    .X(_2948_));
 sky130_fd_sc_hd__xnor2_2 _7332_ (.A(_2943_),
    .B(_2948_),
    .Y(_2949_));
 sky130_fd_sc_hd__and3_1 _7333_ (.A(_3133_),
    .B(_0689_),
    .C(_2789_),
    .X(_2950_));
 sky130_fd_sc_hd__a31o_1 _7334_ (.A1(_3134_),
    .A2(_0559_),
    .A3(_0420_),
    .B1(_2950_),
    .X(_2951_));
 sky130_fd_sc_hd__a21bo_1 _7335_ (.A1(_2766_),
    .A2(_2799_),
    .B1_N(_2765_),
    .X(_2952_));
 sky130_fd_sc_hd__nor2_1 _7336_ (.A(_2787_),
    .B(_2791_),
    .Y(_2953_));
 sky130_fd_sc_hd__a21oi_1 _7337_ (.A1(_2786_),
    .A2(_2792_),
    .B1(_2953_),
    .Y(_2954_));
 sky130_fd_sc_hd__xnor2_1 _7338_ (.A(_2952_),
    .B(_2954_),
    .Y(_2955_));
 sky130_fd_sc_hd__xnor2_1 _7339_ (.A(_2951_),
    .B(_2955_),
    .Y(_2956_));
 sky130_fd_sc_hd__nand2_1 _7340_ (.A(_2237_),
    .B(_1170_),
    .Y(_2957_));
 sky130_fd_sc_hd__or2b_1 _7341_ (.A(_2793_),
    .B_N(_2794_),
    .X(_2959_));
 sky130_fd_sc_hd__a21boi_1 _7342_ (.A1(_2785_),
    .A2(_2796_),
    .B1_N(_2959_),
    .Y(_2960_));
 sky130_fd_sc_hd__xnor2_1 _7343_ (.A(_2819_),
    .B(_2960_),
    .Y(_2961_));
 sky130_fd_sc_hd__nand2_1 _7344_ (.A(_3135_),
    .B(_0559_),
    .Y(_2962_));
 sky130_fd_sc_hd__xnor2_1 _7345_ (.A(_2961_),
    .B(_2962_),
    .Y(_2963_));
 sky130_fd_sc_hd__xnor2_1 _7346_ (.A(_2957_),
    .B(_2963_),
    .Y(_2964_));
 sky130_fd_sc_hd__nand2_1 _7347_ (.A(_3134_),
    .B(_0689_),
    .Y(_2965_));
 sky130_fd_sc_hd__nand2_1 _7348_ (.A(_2138_),
    .B(_1448_),
    .Y(_2966_));
 sky130_fd_sc_hd__xnor2_1 _7349_ (.A(_2965_),
    .B(_2966_),
    .Y(_2967_));
 sky130_fd_sc_hd__xnor2_1 _7350_ (.A(_2964_),
    .B(_2967_),
    .Y(_2968_));
 sky130_fd_sc_hd__xnor2_1 _7351_ (.A(_2956_),
    .B(_2968_),
    .Y(_2970_));
 sky130_fd_sc_hd__nand2_1 _7352_ (.A(_3490_),
    .B(_2018_),
    .Y(_2971_));
 sky130_fd_sc_hd__nand2_1 _7353_ (.A(_3591_),
    .B(_2051_),
    .Y(_2972_));
 sky130_fd_sc_hd__xnor2_1 _7354_ (.A(_2971_),
    .B(_2972_),
    .Y(_2973_));
 sky130_fd_sc_hd__xnor2_1 _7355_ (.A(_2970_),
    .B(_2973_),
    .Y(_2974_));
 sky130_fd_sc_hd__a31o_1 _7356_ (.A1(_2903_),
    .A2(_1778_),
    .A3(_2719_),
    .B1(_2717_),
    .X(_2975_));
 sky130_fd_sc_hd__nand2_1 _7357_ (.A(_2710_),
    .B(_2712_),
    .Y(_2976_));
 sky130_fd_sc_hd__nand2_1 _7358_ (.A(_0063_),
    .B(_1821_),
    .Y(_2977_));
 sky130_fd_sc_hd__nand2_1 _7359_ (.A(_3386_),
    .B(_1963_),
    .Y(_2978_));
 sky130_fd_sc_hd__xor2_1 _7360_ (.A(_2977_),
    .B(_2978_),
    .X(_2979_));
 sky130_fd_sc_hd__xnor2_1 _7361_ (.A(_2976_),
    .B(_2979_),
    .Y(_2981_));
 sky130_fd_sc_hd__nand2_1 _7362_ (.A(_0293_),
    .B(_3128_),
    .Y(_2982_));
 sky130_fd_sc_hd__or2b_1 _7363_ (.A(_2725_),
    .B_N(_2737_),
    .X(_2983_));
 sky130_fd_sc_hd__nand2_1 _7364_ (.A(_2182_),
    .B(_1295_),
    .Y(_2984_));
 sky130_fd_sc_hd__o21ai_2 _7365_ (.A1(_2777_),
    .A2(_2778_),
    .B1(_2776_),
    .Y(_2985_));
 sky130_fd_sc_hd__xnor2_2 _7366_ (.A(_2984_),
    .B(_2985_),
    .Y(_2986_));
 sky130_fd_sc_hd__xnor2_1 _7367_ (.A(_2983_),
    .B(_2986_),
    .Y(_2987_));
 sky130_fd_sc_hd__xnor2_1 _7368_ (.A(_2982_),
    .B(_2987_),
    .Y(_2988_));
 sky130_fd_sc_hd__xnor2_1 _7369_ (.A(_2981_),
    .B(_2988_),
    .Y(_2989_));
 sky130_fd_sc_hd__xnor2_1 _7370_ (.A(_2975_),
    .B(_2989_),
    .Y(_2990_));
 sky130_fd_sc_hd__xnor2_1 _7371_ (.A(_2974_),
    .B(_2990_),
    .Y(_2992_));
 sky130_fd_sc_hd__nand2_1 _7372_ (.A(_2754_),
    .B(_2755_),
    .Y(_2993_));
 sky130_fd_sc_hd__o21ai_1 _7373_ (.A1(_2748_),
    .A2(_2756_),
    .B1(_2993_),
    .Y(_2994_));
 sky130_fd_sc_hd__nand2_1 _7374_ (.A(_2739_),
    .B(_2763_),
    .Y(_2995_));
 sky130_fd_sc_hd__nand2_1 _7375_ (.A(_3209_),
    .B(net57),
    .Y(_2996_));
 sky130_fd_sc_hd__nand2_1 _7376_ (.A(_1045_),
    .B(net54),
    .Y(_2997_));
 sky130_fd_sc_hd__xor2_1 _7377_ (.A(_2996_),
    .B(_2997_),
    .X(_2998_));
 sky130_fd_sc_hd__xnor2_1 _7378_ (.A(_2995_),
    .B(_2998_),
    .Y(_2999_));
 sky130_fd_sc_hd__xnor2_1 _7379_ (.A(_2994_),
    .B(_2999_),
    .Y(_3000_));
 sky130_fd_sc_hd__nand2_1 _7380_ (.A(_0571_),
    .B(_3046_),
    .Y(_3001_));
 sky130_fd_sc_hd__nand2_1 _7381_ (.A(_3425_),
    .B(_1942_),
    .Y(_3003_));
 sky130_fd_sc_hd__nand2_1 _7382_ (.A(_3513_),
    .B(_1909_),
    .Y(_3004_));
 sky130_fd_sc_hd__xnor2_1 _7383_ (.A(_3003_),
    .B(_3004_),
    .Y(_3005_));
 sky130_fd_sc_hd__xnor2_1 _7384_ (.A(_3001_),
    .B(_3005_),
    .Y(_3006_));
 sky130_fd_sc_hd__nand2_1 _7385_ (.A(_2903_),
    .B(_1810_),
    .Y(_3007_));
 sky130_fd_sc_hd__nand2_1 _7386_ (.A(_3720_),
    .B(_0862_),
    .Y(_3008_));
 sky130_fd_sc_hd__and2_1 _7387_ (.A(_2728_),
    .B(_2734_),
    .X(_3009_));
 sky130_fd_sc_hd__a21oi_1 _7388_ (.A1(_2727_),
    .A2(_2735_),
    .B1(_3009_),
    .Y(_3010_));
 sky130_fd_sc_hd__xnor2_1 _7389_ (.A(_3008_),
    .B(_3010_),
    .Y(_3011_));
 sky130_fd_sc_hd__xnor2_1 _7390_ (.A(_3007_),
    .B(_3011_),
    .Y(_3012_));
 sky130_fd_sc_hd__nand2_1 _7391_ (.A(_3486_),
    .B(_2007_),
    .Y(_3014_));
 sky130_fd_sc_hd__xnor2_1 _7392_ (.A(_3012_),
    .B(_3014_),
    .Y(_3015_));
 sky130_fd_sc_hd__xnor2_1 _7393_ (.A(_3006_),
    .B(_3015_),
    .Y(_3016_));
 sky130_fd_sc_hd__xnor2_1 _7394_ (.A(_3000_),
    .B(_3016_),
    .Y(_3017_));
 sky130_fd_sc_hd__xnor2_1 _7395_ (.A(_2992_),
    .B(_3017_),
    .Y(_3018_));
 sky130_fd_sc_hd__xnor2_2 _7396_ (.A(_2949_),
    .B(_3018_),
    .Y(_3019_));
 sky130_fd_sc_hd__xnor2_1 _7397_ (.A(_2938_),
    .B(_3019_),
    .Y(_3020_));
 sky130_fd_sc_hd__xnor2_1 _7398_ (.A(_2937_),
    .B(_3020_),
    .Y(_3021_));
 sky130_fd_sc_hd__xnor2_1 _7399_ (.A(_2931_),
    .B(_3021_),
    .Y(_3022_));
 sky130_fd_sc_hd__xnor2_1 _7400_ (.A(_2930_),
    .B(_3022_),
    .Y(_3023_));
 sky130_fd_sc_hd__and2b_1 _7401_ (.A_N(_2836_),
    .B(_2838_),
    .X(_3025_));
 sky130_fd_sc_hd__a31o_1 _7402_ (.A1(_1067_),
    .A2(net54),
    .A3(_2809_),
    .B1(_2808_),
    .X(_3026_));
 sky130_fd_sc_hd__a21oi_1 _7403_ (.A1(_2779_),
    .A2(_2780_),
    .B1(_2782_),
    .Y(_3027_));
 sky130_fd_sc_hd__xnor2_1 _7404_ (.A(_3026_),
    .B(_3027_),
    .Y(_3028_));
 sky130_fd_sc_hd__or2b_1 _7405_ (.A(_2829_),
    .B_N(_2832_),
    .X(_3029_));
 sky130_fd_sc_hd__nand2_1 _7406_ (.A(_2346_),
    .B(_1949_),
    .Y(_3030_));
 sky130_fd_sc_hd__o21ba_1 _7407_ (.A1(_2815_),
    .A2(_2816_),
    .B1_N(_2813_),
    .X(_3031_));
 sky130_fd_sc_hd__a21oi_1 _7408_ (.A1(_2853_),
    .A2(_2855_),
    .B1(_2852_),
    .Y(_3032_));
 sky130_fd_sc_hd__xnor2_1 _7409_ (.A(_3031_),
    .B(_3032_),
    .Y(_3033_));
 sky130_fd_sc_hd__xnor2_1 _7410_ (.A(_3030_),
    .B(_3033_),
    .Y(_3034_));
 sky130_fd_sc_hd__nand2_1 _7411_ (.A(_2412_),
    .B(_1797_),
    .Y(_3036_));
 sky130_fd_sc_hd__xnor2_1 _7412_ (.A(_3034_),
    .B(_3036_),
    .Y(_3037_));
 sky130_fd_sc_hd__xnor2_1 _7413_ (.A(_2857_),
    .B(_3037_),
    .Y(_3038_));
 sky130_fd_sc_hd__xnor2_1 _7414_ (.A(_3029_),
    .B(_3038_),
    .Y(_3039_));
 sky130_fd_sc_hd__xnor2_1 _7415_ (.A(_3028_),
    .B(_3039_),
    .Y(_3040_));
 sky130_fd_sc_hd__xnor2_1 _7416_ (.A(_3025_),
    .B(_3040_),
    .Y(_3041_));
 sky130_fd_sc_hd__xnor2_1 _7417_ (.A(_3023_),
    .B(_3041_),
    .Y(_3042_));
 sky130_fd_sc_hd__a21oi_1 _7418_ (.A1(_2900_),
    .A2(_3042_),
    .B1(_3192_),
    .Y(_3043_));
 sky130_fd_sc_hd__o21ai_1 _7419_ (.A1(_2900_),
    .A2(_3042_),
    .B1(_3043_),
    .Y(_3044_));
 sky130_fd_sc_hd__o311a_1 _7420_ (.A1(_0181_),
    .A2(_2888_),
    .A3(_2889_),
    .B1(_2899_),
    .C1(_3044_),
    .X(_3045_));
 sky130_fd_sc_hd__nand2_2 _7421_ (.A(_2886_),
    .B(_3045_),
    .Y(net93));
 sky130_fd_sc_hd__mux4_1 _7422_ (.A0(_1067_),
    .A1(_1045_),
    .A2(_1034_),
    .A3(_1023_),
    .S0(_0914_),
    .S1(_0958_),
    .X(_3047_));
 sky130_fd_sc_hd__mux4_1 _7423_ (.A0(_3136_),
    .A1(_3140_),
    .A2(_3138_),
    .A3(_3047_),
    .S0(_1723_),
    .S1(_1712_),
    .X(_3048_));
 sky130_fd_sc_hd__a22o_1 _7424_ (.A1(_3162_),
    .A2(_3487_),
    .B1(_3048_),
    .B2(_0838_),
    .X(_3049_));
 sky130_fd_sc_hd__a21o_1 _7425_ (.A1(_3127_),
    .A2(_0703_),
    .B1(_3049_),
    .X(_3050_));
 sky130_fd_sc_hd__nor2_1 _7426_ (.A(_0860_),
    .B(_0712_),
    .Y(_3051_));
 sky130_fd_sc_hd__a22o_1 _7427_ (.A1(_0925_),
    .A2(_1067_),
    .B1(_3209_),
    .B2(_0969_),
    .X(_3052_));
 sky130_fd_sc_hd__and3b_1 _7428_ (.A_N(_1603_),
    .B(_1668_),
    .C(_3052_),
    .X(_3053_));
 sky130_fd_sc_hd__a221o_1 _7429_ (.A1(_0717_),
    .A2(net123),
    .B1(_1187_),
    .B2(_0685_),
    .C1(_3053_),
    .X(_3054_));
 sky130_fd_sc_hd__or2_1 _7430_ (.A(_0455_),
    .B(_0696_),
    .X(_3055_));
 sky130_fd_sc_hd__nand2_1 _7431_ (.A(_0455_),
    .B(_0696_),
    .Y(_3057_));
 sky130_fd_sc_hd__o21ba_1 _7432_ (.A1(_0717_),
    .A2(_1209_),
    .B1_N(_1220_),
    .X(_3058_));
 sky130_fd_sc_hd__xor2_1 _7433_ (.A(_0455_),
    .B(_0510_),
    .X(_3059_));
 sky130_fd_sc_hd__a2bb2o_1 _7434_ (.A1_N(_0685_),
    .A2_N(_3058_),
    .B1(_3059_),
    .B2(_0652_),
    .X(_3060_));
 sky130_fd_sc_hd__a31o_1 _7435_ (.A1(_3055_),
    .A2(_2980_),
    .A3(_3057_),
    .B1(_3060_),
    .X(_3061_));
 sky130_fd_sc_hd__a2111o_4 _7436_ (.A1(_3587_),
    .A2(_3050_),
    .B1(_3051_),
    .C1(_3054_),
    .D1(_3061_),
    .X(net80));
 sky130_fd_sc_hd__nor2_1 _7437_ (.A(_2672_),
    .B(_2697_),
    .Y(_3062_));
 sky130_fd_sc_hd__o21a_1 _7438_ (.A1(_2672_),
    .A2(_2677_),
    .B1(_2701_),
    .X(_3063_));
 sky130_fd_sc_hd__o211ai_1 _7439_ (.A1(_2697_),
    .A2(_3063_),
    .B1(_2887_),
    .C1(_2883_),
    .Y(_3064_));
 sky130_fd_sc_hd__a31o_1 _7440_ (.A1(_2303_),
    .A2(_2309_),
    .A3(_3062_),
    .B1(_3064_),
    .X(_3065_));
 sky130_fd_sc_hd__or2b_1 _7441_ (.A(net57),
    .B_N(_0571_),
    .X(_3067_));
 sky130_fd_sc_hd__or4b_1 _7442_ (.A(_1165_),
    .B(_0783_),
    .C(_1144_),
    .D_N(_1154_),
    .X(_3068_));
 sky130_fd_sc_hd__a21o_1 _7443_ (.A1(_3065_),
    .A2(_3067_),
    .B1(_3068_),
    .X(_3069_));
 sky130_fd_sc_hd__a21o_1 _7444_ (.A1(_0863_),
    .A2(_1067_),
    .B1(_3211_),
    .X(_3070_));
 sky130_fd_sc_hd__mux2_1 _7445_ (.A0(_1045_),
    .A1(_1034_),
    .S(_0925_),
    .X(_3071_));
 sky130_fd_sc_hd__mux4_1 _7446_ (.A0(_2357_),
    .A1(_3070_),
    .A2(_2467_),
    .A3(_3071_),
    .S0(_0866_),
    .S1(_0864_),
    .X(_3072_));
 sky130_fd_sc_hd__mux4_1 _7447_ (.A0(_3400_),
    .A1(_3403_),
    .A2(_3072_),
    .A3(_3401_),
    .S0(_0861_),
    .S1(_0867_),
    .X(_3073_));
 sky130_fd_sc_hd__nand2_2 _7448_ (.A(_3587_),
    .B(_3073_),
    .Y(_3074_));
 sky130_fd_sc_hd__and2_1 _7449_ (.A(_0510_),
    .B(_3210_),
    .X(_3075_));
 sky130_fd_sc_hd__o22a_1 _7450_ (.A1(_3305_),
    .A2(_0696_),
    .B1(_0438_),
    .B2(_3075_),
    .X(_3076_));
 sky130_fd_sc_hd__o32a_1 _7451_ (.A1(_0863_),
    .A2(_3209_),
    .A3(_0855_),
    .B1(_3076_),
    .B2(_1277_),
    .X(_3078_));
 sky130_fd_sc_hd__inv_2 _7452_ (.A(_3078_),
    .Y(_3079_));
 sky130_fd_sc_hd__o22a_1 _7453_ (.A1(_0696_),
    .A2(_0309_),
    .B1(_3075_),
    .B2(_0641_),
    .X(_3080_));
 sky130_fd_sc_hd__o311a_1 _7454_ (.A1(_0860_),
    .A2(_3210_),
    .A3(_0196_),
    .B1(_3079_),
    .C1(_3080_),
    .X(_3081_));
 sky130_fd_sc_hd__nand3_4 _7455_ (.A(_3069_),
    .B(_3074_),
    .C(_3081_),
    .Y(net69));
 sky130_fd_sc_hd__mux4_1 _7456_ (.A0(_1034_),
    .A1(_2346_),
    .A2(_1023_),
    .A3(_2412_),
    .S0(_0947_),
    .S1(_0914_),
    .X(_3082_));
 sky130_fd_sc_hd__mux4_1 _7457_ (.A0(_3298_),
    .A1(_3300_),
    .A2(_3299_),
    .A3(_3082_),
    .S0(_0587_),
    .S1(_1712_),
    .X(_3083_));
 sky130_fd_sc_hd__mux2_1 _7458_ (.A0(_0885_),
    .A1(_3083_),
    .S(_0838_),
    .X(_3084_));
 sky130_fd_sc_hd__a41o_1 _7459_ (.A1(_3127_),
    .A2(net25),
    .A3(_0783_),
    .A4(_1734_),
    .B1(_3084_),
    .X(_3085_));
 sky130_fd_sc_hd__o21ai_1 _7460_ (.A1(_1613_),
    .A2(_1635_),
    .B1(_1668_),
    .Y(_3086_));
 sky130_fd_sc_hd__a21oi_1 _7461_ (.A1(_0237_),
    .A2(_3158_),
    .B1(_1220_),
    .Y(_3088_));
 sky130_fd_sc_hd__o22a_1 _7462_ (.A1(_0860_),
    .A2(_0869_),
    .B1(_3088_),
    .B2(_0674_),
    .X(_3089_));
 sky130_fd_sc_hd__o221a_1 _7463_ (.A1(_0237_),
    .A2(_0309_),
    .B1(_3712_),
    .B2(_0248_),
    .C1(_3089_),
    .X(_3090_));
 sky130_fd_sc_hd__and2_1 _7464_ (.A(_0259_),
    .B(_0576_),
    .X(_3091_));
 sky130_fd_sc_hd__nor2_1 _7465_ (.A(_0259_),
    .B(_0576_),
    .Y(_3092_));
 sky130_fd_sc_hd__xnor2_1 _7466_ (.A(_0259_),
    .B(_0761_),
    .Y(_3093_));
 sky130_fd_sc_hd__o32a_1 _7467_ (.A1(_3091_),
    .A2(_3265_),
    .A3(_3092_),
    .B1(_3093_),
    .B2(_3595_),
    .X(_3094_));
 sky130_fd_sc_hd__o211a_1 _7468_ (.A1(_1646_),
    .A2(_3086_),
    .B1(_3090_),
    .C1(_3094_),
    .X(_3095_));
 sky130_fd_sc_hd__a21bo_1 _7469_ (.A1(_1701_),
    .A2(_3085_),
    .B1_N(_3095_),
    .X(_3096_));
 sky130_fd_sc_hd__buf_2 _7470_ (.A(_3096_),
    .X(net94));
 sky130_fd_sc_hd__mux4_1 _7471_ (.A0(_2467_),
    .A1(_3071_),
    .A2(_2193_),
    .A3(_2357_),
    .S0(_3077_),
    .S1(_0969_),
    .X(_3098_));
 sky130_fd_sc_hd__mux4_1 _7472_ (.A0(_3581_),
    .A1(_3584_),
    .A2(_3098_),
    .A3(_3582_),
    .S0(_0063_),
    .S1(_3301_),
    .X(_3099_));
 sky130_fd_sc_hd__nand2_1 _7473_ (.A(_0379_),
    .B(_0728_),
    .Y(_3100_));
 sky130_fd_sc_hd__or2_1 _7474_ (.A(_0379_),
    .B(_0728_),
    .X(_3101_));
 sky130_fd_sc_hd__a21oi_1 _7475_ (.A1(_0379_),
    .A2(_0543_),
    .B1(_3265_),
    .Y(_3102_));
 sky130_fd_sc_hd__o21a_1 _7476_ (.A1(_0379_),
    .A2(_0543_),
    .B1(_3102_),
    .X(_3103_));
 sky130_fd_sc_hd__a31o_1 _7477_ (.A1(_2980_),
    .A2(_3100_),
    .A3(_3101_),
    .B1(_3103_),
    .X(_3104_));
 sky130_fd_sc_hd__a31o_1 _7478_ (.A1(_3490_),
    .A2(_3591_),
    .A3(_3162_),
    .B1(_3104_),
    .X(_3105_));
 sky130_fd_sc_hd__o21ai_1 _7479_ (.A1(_1592_),
    .A2(_1603_),
    .B1(_1668_),
    .Y(_3106_));
 sky130_fd_sc_hd__a21oi_1 _7480_ (.A1(_0750_),
    .A2(_3158_),
    .B1(_3204_),
    .Y(_3107_));
 sky130_fd_sc_hd__a22oi_1 _7481_ (.A1(_0270_),
    .A2(net123),
    .B1(_1187_),
    .B2(_0368_),
    .Y(_3109_));
 sky130_fd_sc_hd__o221a_1 _7482_ (.A1(_0860_),
    .A2(_0850_),
    .B1(_3107_),
    .B2(_0368_),
    .C1(_3109_),
    .X(_3110_));
 sky130_fd_sc_hd__o21ai_1 _7483_ (.A1(_1613_),
    .A2(_3106_),
    .B1(_3110_),
    .Y(_3111_));
 sky130_fd_sc_hd__a211o_1 _7484_ (.A1(_3587_),
    .A2(_3099_),
    .B1(_3105_),
    .C1(_3111_),
    .X(net91));
 sky130_fd_sc_hd__or3_1 _7485_ (.A(net86),
    .B(net87),
    .C(net89),
    .X(_3112_));
 sky130_fd_sc_hd__or4_1 _7486_ (.A(net95),
    .B(net80),
    .C(net94),
    .D(net91),
    .X(_3113_));
 sky130_fd_sc_hd__or4_1 _7487_ (.A(net96),
    .B(net97),
    .C(net98),
    .D(_3113_),
    .X(_3114_));
 sky130_fd_sc_hd__or3_1 _7488_ (.A(net99),
    .B(net100),
    .C(_3114_),
    .X(_3115_));
 sky130_fd_sc_hd__or3_1 _7489_ (.A(net70),
    .B(net71),
    .C(_3115_),
    .X(_3116_));
 sky130_fd_sc_hd__or4_1 _7490_ (.A(net72),
    .B(net73),
    .C(net74),
    .D(_3116_),
    .X(_3117_));
 sky130_fd_sc_hd__or4_2 _7491_ (.A(net75),
    .B(net76),
    .C(net77),
    .D(_3117_),
    .X(_3119_));
 sky130_fd_sc_hd__nor4_1 _7492_ (.A(net78),
    .B(net79),
    .C(net81),
    .D(_3119_),
    .Y(_3120_));
 sky130_fd_sc_hd__and4b_1 _7493_ (.A_N(net85),
    .B(_3069_),
    .C(_3074_),
    .D(_3081_),
    .X(_3121_));
 sky130_fd_sc_hd__and4bb_1 _7494_ (.A_N(net82),
    .B_N(net83),
    .C(_3120_),
    .D(_3121_),
    .X(_3122_));
 sky130_fd_sc_hd__nor4b_1 _7495_ (.A(net88),
    .B(_2669_),
    .C(_2676_),
    .D_N(_2692_),
    .Y(_3123_));
 sky130_fd_sc_hd__and4bb_1 _7496_ (.A_N(net84),
    .B_N(_3112_),
    .C(_3122_),
    .D(_3123_),
    .X(_3124_));
 sky130_fd_sc_hd__and4b_2 _7497_ (.A_N(net92),
    .B(_2886_),
    .C(_3045_),
    .D(_3124_),
    .X(_3125_));
 sky130_fd_sc_hd__buf_6 _7498_ (.A(_3125_),
    .X(net101));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__buf_4 input1 (.A(A[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(A[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input3 (.A(A[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(A[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(A[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(A[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(A[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(A[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input9 (.A(A[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_4 input10 (.A(A[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_8 input11 (.A(A[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_6 input12 (.A(A[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_4 input13 (.A(A[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(A[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input15 (.A(A[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_4 input16 (.A(A[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_4 input17 (.A(A[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 input18 (.A(A[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input19 (.A(A[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_4 input20 (.A(A[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_4 input21 (.A(A[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(A[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_4 input23 (.A(A[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(A[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_4 input25 (.A(A[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 input26 (.A(A[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_6 input27 (.A(A[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_4 input28 (.A(A[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_4 input29 (.A(A[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 input30 (.A(A[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_8 input31 (.A(A[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_4 input32 (.A(A[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_6 input33 (.A(B[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(B[10]),
    .X(net34));
 sky130_fd_sc_hd__buf_2 input35 (.A(B[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 input36 (.A(B[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_2 input37 (.A(B[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_4 input38 (.A(B[14]),
    .X(net38));
 sky130_fd_sc_hd__buf_2 input39 (.A(B[15]),
    .X(net39));
 sky130_fd_sc_hd__buf_2 input40 (.A(B[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 input41 (.A(B[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(B[18]),
    .X(net42));
 sky130_fd_sc_hd__buf_2 input43 (.A(B[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_4 input44 (.A(B[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 input45 (.A(B[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 input46 (.A(B[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 input47 (.A(B[22]),
    .X(net47));
 sky130_fd_sc_hd__buf_4 input48 (.A(B[23]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(B[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 input50 (.A(B[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_4 input51 (.A(B[26]),
    .X(net51));
 sky130_fd_sc_hd__buf_2 input52 (.A(B[27]),
    .X(net52));
 sky130_fd_sc_hd__buf_2 input53 (.A(B[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_4 input54 (.A(B[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_2 input55 (.A(B[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_8 input56 (.A(B[30]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 input57 (.A(B[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_6 input58 (.A(B[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_4 input59 (.A(B[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_8 input60 (.A(B[5]),
    .X(net60));
 sky130_fd_sc_hd__buf_8 input61 (.A(B[6]),
    .X(net61));
 sky130_fd_sc_hd__buf_6 input62 (.A(B[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_2 input63 (.A(B[8]),
    .X(net63));
 sky130_fd_sc_hd__buf_4 input64 (.A(B[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_4 input65 (.A(control[0]),
    .X(net65));
 sky130_fd_sc_hd__buf_2 input66 (.A(control[1]),
    .X(net66));
 sky130_fd_sc_hd__buf_4 input67 (.A(control[2]),
    .X(net67));
 sky130_fd_sc_hd__buf_2 input68 (.A(control[3]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net69),
    .X(result[0]));
 sky130_fd_sc_hd__clkbuf_4 output70 (.A(net70),
    .X(result[10]));
 sky130_fd_sc_hd__clkbuf_4 output71 (.A(net71),
    .X(result[11]));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net72),
    .X(result[12]));
 sky130_fd_sc_hd__clkbuf_4 output73 (.A(net73),
    .X(result[13]));
 sky130_fd_sc_hd__clkbuf_4 output74 (.A(net74),
    .X(result[14]));
 sky130_fd_sc_hd__clkbuf_4 output75 (.A(net75),
    .X(result[15]));
 sky130_fd_sc_hd__clkbuf_4 output76 (.A(net76),
    .X(result[16]));
 sky130_fd_sc_hd__clkbuf_4 output77 (.A(net77),
    .X(result[17]));
 sky130_fd_sc_hd__clkbuf_4 output78 (.A(net78),
    .X(result[18]));
 sky130_fd_sc_hd__clkbuf_4 output79 (.A(net79),
    .X(result[19]));
 sky130_fd_sc_hd__clkbuf_4 output80 (.A(net80),
    .X(result[1]));
 sky130_fd_sc_hd__clkbuf_4 output81 (.A(net81),
    .X(result[20]));
 sky130_fd_sc_hd__clkbuf_4 output82 (.A(net82),
    .X(result[21]));
 sky130_fd_sc_hd__clkbuf_4 output83 (.A(net83),
    .X(result[22]));
 sky130_fd_sc_hd__clkbuf_4 output84 (.A(net84),
    .X(result[23]));
 sky130_fd_sc_hd__clkbuf_4 output85 (.A(net167),
    .X(result[24]));
 sky130_fd_sc_hd__clkbuf_4 output86 (.A(net86),
    .X(result[25]));
 sky130_fd_sc_hd__clkbuf_4 output87 (.A(net166),
    .X(result[26]));
 sky130_fd_sc_hd__clkbuf_4 output88 (.A(net88),
    .X(result[27]));
 sky130_fd_sc_hd__clkbuf_4 output89 (.A(net89),
    .X(result[28]));
 sky130_fd_sc_hd__clkbuf_4 output90 (.A(net90),
    .X(result[29]));
 sky130_fd_sc_hd__clkbuf_4 output91 (.A(net91),
    .X(result[2]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(result[30]));
 sky130_fd_sc_hd__clkbuf_4 output93 (.A(net93),
    .X(result[31]));
 sky130_fd_sc_hd__clkbuf_4 output94 (.A(net94),
    .X(result[3]));
 sky130_fd_sc_hd__clkbuf_4 output95 (.A(net165),
    .X(result[4]));
 sky130_fd_sc_hd__clkbuf_4 output96 (.A(net96),
    .X(result[5]));
 sky130_fd_sc_hd__clkbuf_4 output97 (.A(net97),
    .X(result[6]));
 sky130_fd_sc_hd__clkbuf_4 output98 (.A(net98),
    .X(result[7]));
 sky130_fd_sc_hd__clkbuf_4 output99 (.A(net99),
    .X(result[8]));
 sky130_fd_sc_hd__clkbuf_4 output100 (.A(net100),
    .X(result[9]));
 sky130_fd_sc_hd__buf_6 output101 (.A(net101),
    .X(zero_flag));
 sky130_fd_sc_hd__buf_1 max_cap102 (.A(_2849_),
    .X(net102));
 sky130_fd_sc_hd__buf_1 max_cap103 (.A(_1989_),
    .X(net103));
 sky130_fd_sc_hd__buf_1 wire104 (.A(net200),
    .X(net104));
 sky130_fd_sc_hd__buf_1 max_cap105 (.A(_1814_),
    .X(net105));
 sky130_fd_sc_hd__buf_1 wire106 (.A(_0986_),
    .X(net106));
 sky130_fd_sc_hd__buf_1 max_cap107 (.A(_1191_),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 max_cap108 (.A(_1737_),
    .X(net108));
 sky130_fd_sc_hd__buf_1 max_cap109 (.A(_1420_),
    .X(net109));
 sky130_fd_sc_hd__buf_1 max_cap110 (.A(net111),
    .X(net110));
 sky130_fd_sc_hd__buf_1 wire111 (.A(_1068_),
    .X(net111));
 sky130_fd_sc_hd__buf_1 max_cap112 (.A(_0803_),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 max_cap113 (.A(_0648_),
    .X(net113));
 sky130_fd_sc_hd__buf_1 max_cap114 (.A(_0398_),
    .X(net114));
 sky130_fd_sc_hd__buf_1 max_cap115 (.A(net202),
    .X(net115));
 sky130_fd_sc_hd__buf_1 max_cap116 (.A(_0155_),
    .X(net116));
 sky130_fd_sc_hd__buf_1 max_cap117 (.A(_2186_),
    .X(net117));
 sky130_fd_sc_hd__buf_1 max_cap118 (.A(_1088_),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 max_cap119 (.A(_0979_),
    .X(net119));
 sky130_fd_sc_hd__buf_1 max_cap120 (.A(_1904_),
    .X(net120));
 sky130_fd_sc_hd__buf_1 max_cap121 (.A(_1543_),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_2 max_cap122 (.A(_3370_),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 max_cap123 (.A(_1176_),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 max_cap124 (.A(_3158_),
    .X(net124));
 sky130_fd_sc_hd__buf_1 rebuffer1 (.A(_0526_),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 rebuffer2 (.A(_3682_),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 rebuffer3 (.A(net126),
    .X(net127));
 sky130_fd_sc_hd__buf_1 rebuffer4 (.A(_1121_),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 rebuffer5 (.A(net153),
    .X(net129));
 sky130_fd_sc_hd__buf_1 rebuffer6 (.A(_0984_),
    .X(net130));
 sky130_fd_sc_hd__buf_1 rebuffer7 (.A(_3529_),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 rebuffer8 (.A(_0993_),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 rebuffer9 (.A(net132),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 rebuffer10 (.A(_1135_),
    .X(net134));
 sky130_fd_sc_hd__buf_1 rebuffer11 (.A(_0650_),
    .X(net135));
 sky130_fd_sc_hd__buf_1 rebuffer12 (.A(_1126_),
    .X(net136));
 sky130_fd_sc_hd__buf_6 rebuffer13 (.A(_1126_),
    .X(net137));
 sky130_fd_sc_hd__buf_1 rebuffer14 (.A(_3666_),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 rebuffer15 (.A(net138),
    .X(net139));
 sky130_fd_sc_hd__buf_1 rebuffer16 (.A(_0679_),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 rebuffer17 (.A(net140),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 rebuffer18 (.A(_0083_),
    .X(net142));
 sky130_fd_sc_hd__buf_1 rebuffer19 (.A(_2047_),
    .X(net143));
 sky130_fd_sc_hd__buf_6 rebuffer20 (.A(_3556_),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 rebuffer21 (.A(_3257_),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 rebuffer22 (.A(_3257_),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 rebuffer23 (.A(_3257_),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 rebuffer24 (.A(_3674_),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer25 (.A(net148),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 rebuffer26 (.A(net148),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 rebuffer27 (.A(net150),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 rebuffer28 (.A(_2147_),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 rebuffer29 (.A(_1619_),
    .X(net153));
 sky130_fd_sc_hd__buf_1 rebuffer30 (.A(_1422_),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 rebuffer31 (.A(_3628_),
    .X(net155));
 sky130_fd_sc_hd__buf_1 rebuffer32 (.A(_0271_),
    .X(net156));
 sky130_fd_sc_hd__buf_1 rebuffer33 (.A(_2098_),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 rebuffer34 (.A(_2098_),
    .X(net158));
 sky130_fd_sc_hd__buf_1 rebuffer35 (.A(_3255_),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 rebuffer36 (.A(net159),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 rebuffer37 (.A(_1134_),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_2 split38 (.A(_3270_),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 split39 (.A(_0412_),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 rebuffer40 (.A(_0552_),
    .X(net164));
 sky130_fd_sc_hd__buf_2 rebuffer41 (.A(net95),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_4 rebuffer42 (.A(net87),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_4 rebuffer43 (.A(net85),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 rebuffer44 (.A(_2493_),
    .X(net168));
 sky130_fd_sc_hd__buf_1 rebuffer45 (.A(_2096_),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_1 rebuffer46 (.A(_2096_),
    .X(net170));
 sky130_fd_sc_hd__buf_1 rebuffer47 (.A(_2101_),
    .X(net171));
 sky130_fd_sc_hd__buf_1 rebuffer48 (.A(net115),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer49 (.A(_0396_),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 rebuffer50 (.A(_1921_),
    .X(net174));
 sky130_fd_sc_hd__buf_1 rebuffer51 (.A(_1921_),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 rebuffer52 (.A(_3259_),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 rebuffer53 (.A(_2111_),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_2 split54 (.A(_3176_),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 rebuffer55 (.A(_0405_),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_1 rebuffer56 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_1 rebuffer57 (.A(_0408_),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 rebuffer58 (.A(_2094_),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 rebuffer59 (.A(_3372_),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 rebuffer60 (.A(_3371_),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 rebuffer61 (.A(_1915_),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 rebuffer62 (.A(_3374_),
    .X(net186));
 sky130_fd_sc_hd__buf_1 rebuffer63 (.A(_1086_),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 rebuffer64 (.A(_3379_),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer65 (.A(_2025_),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 rebuffer66 (.A(_0267_),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_2 split67 (.A(_0030_),
    .X(net191));
 sky130_fd_sc_hd__buf_1 rebuffer68 (.A(_3334_),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer69 (.A(_3233_),
    .X(net193));
 sky130_fd_sc_hd__buf_6 split70 (.A(_0074_),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_1 rebuffer71 (.A(_3178_),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_1 rebuffer72 (.A(_3376_),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_1 max_cap1 (.A(_2849_),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_1 max_cap2 (.A(_1324_),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 max_cap3 (.A(_1158_),
    .X(net199));
 sky130_fd_sc_hd__buf_1 wire4 (.A(_2052_),
    .X(net200));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_cap5 (.A(_1737_),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_1 max_cap6 (.A(_0398_),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 max_cap7 (.A(_1420_),
    .X(net203));
endmodule
